Standard cell Simulation
* takes 3:47 to run

.include "/home/matt/work/asic-workshop/shuttle5/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt.spice"
* include this one, so that don't need to extract models with magic
.include "/home/matt/work/asic-workshop/shuttle5/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice"
* now we can just use the spice file generated in the openlane run
.include "instrumented_adder.spice"

* instantiate the spice model
* Xpoc  chain clk outputs[0] outputs[1] outputs[2] outputs[3] reset VPWR VGND instrumented_adder
Xpoc b[0] b[1] b[2] b[3] b[4] b[5] b[6] b[7] bypass chain clk
+ extra_inverter reset ring_osc_counter_out[0] ring_osc_counter_out[1] ring_osc_counter_out[2]
+ ring_osc_counter_out[3] ring_osc_counter_out[4] ring_osc_counter_out[5] ring_osc_counter_out[6]
+ ring_osc_counter_out[7] run time_count_overflow VPWR VGND instrumented_adder

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8
Vbypass bypass VGND 0
Vextra_inverter extra_inverter VGND 1.8
Vrun run VGND 1.8

* b input
Vb0 b[0] VGND 1.8
Vb1 b[1] VGND 0
Vb2 b[2] VGND 0
Vb3 b[3] VGND 0
Vb4 b[4] VGND 0
Vb5 b[5] VGND 0
Vb6 b[6] VGND 0
Vb7 b[7] VGND 0

* create a clock, 4ns period
* initial v, pulse v, delay, rise, fall, pulse w, period
Vclk clk VGND pulse(0 1.8 1n 10p 10p 2n 4n)

* create reset
* start high, for 2ns, rest of the time off
Vreset reset VGND pulse(0 1.8 0n 10p 10p 2n 20n)

* setup the transient analysis
.tran 10p 10n 0

.control
run
set color0 = white
set color1 = black
plot reset, clk, chain, time_count_overflow
.endc

.end
