Standard cell Simulation

.include "/home/matt/work/asic-workshop/shuttle5/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt.spice"
.include "instrumented_adder.spice"

* instantiate the spice model
Xpoc  chain clk outputs[0] outputs[1] outputs[2] outputs[3] reset VPWR VGND instrumented_adder

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create a clock, 4ns period
* initial v, pulse v, delay, rise, fall, pulse w, period
Vclk clk VGND pulse(0 1.8 1n 10p 10p 2n 4n)

* create reset
* start high, for 2ns, rest of the time off
Vreset reset VGND pulse(0 1.8 0n 10p 10p 2n 20n)

* setup the transient analysis
.tran 50p 10n 0

.control
run
set color0 = white
set color1 = black
plot reset, clk, chain
.endc

.end
