latest_run/results/finishing/instrumented_adder.spice