adder kogge_stone

.include "/home/matt/work/asic-workshop/shuttle5/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt.spice"
* include this one, so that don't need to extract models with magic
.include "/home/matt/work/asic-workshop/shuttle5/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice"
* now we can just use the spice file generated in the openlane run
.include "instrumented_adder.spice.kogge_stone"

* instantiate the spice model
Xpoc a_input[0] a_input[1] a_input[2] a_input[3] a_input[4]
+ a_input[5] a_input[6] a_input[7] a_input_ext_bit_b[0] a_input_ext_bit_b[1] a_input_ext_bit_b[2]
+ a_input_ext_bit_b[3] a_input_ext_bit_b[4] a_input_ext_bit_b[5] a_input_ext_bit_b[6]
+ a_input_ext_bit_b[7] a_input_ring_bit_b[0] a_input_ring_bit_b[1] a_input_ring_bit_b[2]
+ a_input_ring_bit_b[3] a_input_ring_bit_b[4] a_input_ring_bit_b[5] a_input_ring_bit_b[6]
+ a_input_ring_bit_b[7] b_input[0] b_input[1] b_input[2] b_input[3] b_input[4] b_input[5]
+ b_input[6] b_input[7] bypass_b clk control_b counter_enable counter_load done extra_inverter
+ integration_time[0] integration_time[10] integration_time[11] integration_time[12]
+ integration_time[13] integration_time[14] integration_time[15] integration_time[16]
+ integration_time[17] integration_time[18] integration_time[19] integration_time[1]
+ integration_time[20] integration_time[21] integration_time[22] integration_time[23]
+ integration_time[24] integration_time[25] integration_time[26] integration_time[27]
+ integration_time[28] integration_time[29] integration_time[2] integration_time[30]
+ integration_time[31] integration_time[3] integration_time[4] integration_time[5]
+ integration_time[6] integration_time[7] integration_time[8] integration_time[9]
+ reset ring_osc_counter_out[0] ring_osc_counter_out[10] ring_osc_counter_out[11]
+ ring_osc_counter_out[12] ring_osc_counter_out[13] ring_osc_counter_out[14] ring_osc_counter_out[15]
+ ring_osc_counter_out[16] ring_osc_counter_out[17] ring_osc_counter_out[18] ring_osc_counter_out[19]
+ ring_osc_counter_out[1] ring_osc_counter_out[20] ring_osc_counter_out[21] ring_osc_counter_out[22]
+ ring_osc_counter_out[23] ring_osc_counter_out[24] ring_osc_counter_out[25] ring_osc_counter_out[26]
+ ring_osc_counter_out[27] ring_osc_counter_out[28] ring_osc_counter_out[29] ring_osc_counter_out[2]
+ ring_osc_counter_out[30] ring_osc_counter_out[31] ring_osc_counter_out[3] ring_osc_counter_out[4]
+ ring_osc_counter_out[5] ring_osc_counter_out[6] ring_osc_counter_out[7] ring_osc_counter_out[8]
+ ring_osc_counter_out[9] ring_osc_out s_output_bit_b[0] s_output_bit_b[1] s_output_bit_b[2]
+ s_output_bit_b[3] s_output_bit_b[4] s_output_bit_b[5] s_output_bit_b[6] s_output_bit_b[7]
+ stop_b sum_out[0] sum_out[1] sum_out[2] sum_out[3] sum_out[4] sum_out[5] sum_out[6]
+ sum_out[7] VPWR VGND instrumented_adder

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8
Vreset reset VGND 1.8
Vbypass_b bypass_b VGND 1.8
Vcontrol_b control_b VGND 1.8
Vextra_inverter extra_inverter VGND 1.8

* a input
Va0 a_input[0] VGND 0
Va1 a_input[1] VGND 0
Va2 a_input[2] VGND 0
Va3 a_input[3] VGND 0
Va4 a_input[4] VGND 0
Va5 a_input[5] VGND 0
Va6 a_input[6] VGND 0
Va7 a_input[7] VGND 0

* b input
Vb0 b_input[0] VGND 0
Vb1 b_input[1] VGND 0
Vb2 b_input[2] VGND 0
Vb3 b_input[3] VGND 0
Vb4 b_input[4] VGND 0
Vb5 b_input[5] VGND 0
Vb6 b_input[6] VGND 0
Vb7 b_input[7] VGND 0

* sum output bit enable
Vob0 s_output_bit_b[0] VGND 1.8
Vob1 s_output_bit_b[1] VGND 1.8
Vob2 s_output_bit_b[2] VGND 1.8
Vob3 s_output_bit_b[3] VGND 1.8
Vob4 s_output_bit_b[4] VGND 1.8
Vob5 s_output_bit_b[5] VGND 1.8
Vob6 s_output_bit_b[6] VGND 1.8
Vob7 s_output_bit_b[7] VGND 0

* a input ring bit select
Vrb0 a_input_ring_bit_b[0] VGND 1.8
Vrb1 a_input_ring_bit_b[1] VGND 1.8
Vrb2 a_input_ring_bit_b[2] VGND 1.8
Vrb3 a_input_ring_bit_b[3] VGND 1.8
Vrb4 a_input_ring_bit_b[4] VGND 1.8
Vrb5 a_input_ring_bit_b[5] VGND 1.8
Vrb6 a_input_ring_bit_b[6] VGND 1.8
Vrb7 a_input_ring_bit_b[7] VGND 0

* a input external bit select
Veb0 a_input_ext_bit_b[0] VGND 0
Veb1 a_input_ext_bit_b[1] VGND 0
Veb2 a_input_ext_bit_b[2] VGND 0
Veb3 a_input_ext_bit_b[3] VGND 0
Veb4 a_input_ext_bit_b[4] VGND 0
Veb5 a_input_ext_bit_b[5] VGND 0
Veb6 a_input_ext_bit_b[6] VGND 0
Veb7 a_input_ext_bit_b[7] VGND 1.8

* create a clock, 4ns period
* initial v, pulse v, delay, rise, fall, pulse w, period
Vclk clk VGND pulse(0 1.8 2n 10p 10p 2n 4n)

* create run signal
Vstop_b stop_b VGND     pulse(0 1.8 2n 10p 10p 200n 300n)

* setup the transient analysis
.tran 10p 8n 0 uic
.meas tran loop_period trig v(ring_osc_out) val='1.4' rise=2 targ v(ring_osc_out) val='1.4' rise=3
.meas tran rise_time   trig v(ring_osc_out) val='0.2' rise=1 targ v(ring_osc_out) val='1.6' rise=2

.control
run
set color0 = white
set color1 = black
plot stop_b, ring_osc_out
.endc

.end
