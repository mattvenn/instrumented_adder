Standard cell Simulation

.include "/home/matt/work/asic-workshop/shuttle5/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt.spice"
* include this one, so that don't need to extract models with magic
.include "/home/matt/work/asic-workshop/shuttle5/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice"
* now we can just use the spice file generated in the openlane run
.include "instrumented_adder.spice"

* instantiate the spice model
* Xpoc  chain clk outputs[0] outputs[1] outputs[2] outputs[3] reset VPWR VGND instrumented_adder
Xpoc b[0] b[1] b[2] b[3] b[4] b[5] b[6] b[7] bypass chain clk
+ counter_end[0] counter_end[1] counter_end[2] counter_end[3]
+ counter_end[4] counter_end[5] counter_end[6] counter_end[7]
+ counter_out[0] counter_out[1] counter_out[2] counter_out[3]
+ counter_out[4] counter_out[5] counter_out[6] counter_out[7]
+ extra_inverter reset ring_osc_counter_out[0] ring_osc_counter_out[1] ring_osc_counter_out[2]
+ ring_osc_counter_out[3] ring_osc_counter_out[4] ring_osc_counter_out[5] ring_osc_counter_out[6]
+ ring_osc_counter_out[7] run time_count_overflow VPWR VGND instrumented_adder

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8
Vbypass bypass VGND 0
Vextra_inverter extra_inverter VGND 1.8
Vrun run VGND 1.8

* b input
Vb0 b[0] VGND 1.8
Vb1 b[1] VGND 0
Vb2 b[2] VGND 0
Vb3 b[3] VGND 0
Vb4 b[4] VGND 0
Vb5 b[5] VGND 0
Vb6 b[6] VGND 0
Vb7 b[7] VGND 0

* count end input: set to 8
Vc0 counter_end[0] VGND 0
Vc1 counter_end[1] VGND 0
Vc2 counter_end[2] VGND 0
Vc3 counter_end[3] VGND 1.8
Vc4 counter_end[4] VGND 0
Vc5 counter_end[5] VGND 0
Vc6 counter_end[6] VGND 0
Vc7 counter_end[7] VGND 0


* create a clock, 4ns period 
* initial v, pulse v, delay, rise, fall, pulse w, period
Vclk clk VGND pulse(0 1.8 2n 10p 10p 2n 4n)

* create reset
* start high, for 100ns, rest of the time off
Vreset reset VGND pulse(0 1.8 1n 10p 10p 4n 200n)

* create run signal
Vrun run VGND     pulse(0 1.8 6n 10p 10p 200n 300n)

* setup the transient analysis
.tran 10p 12n 0 uic
.meas tran loop_period trig v(chain) val='0.9' rise=2 targ v(chain) val='0.9' rise=3
*.meas tran overflow        trig v(run)   val='0.5*Vdd' rise=1 targ v(time_count_overflow)  val='0.5*Vdd' rise=1

.control
run
set color0 = white
set color1 = black
plot reset, chain, run
.endc

.end
