
module ripple_carry(

	input [31:0] a_in,
	input [31:0] b_in,
	output [31:0] sum
	);

// adder_forest tree_31
	wire n124_tree_31, n125_tree_31, n126_tree_31, n127_tree_31, n128_tree_31, n129_tree_31, n130_tree_31, n131_tree_31, n132_tree_31, n133_tree_31, n134_tree_31, n135_tree_31, n136_tree_31, n137_tree_31, n138_tree_31, n139_tree_31, n140_tree_31, n141_tree_31, n142_tree_31, n143_tree_31, n144_tree_31, n145_tree_31, n146_tree_31, n147_tree_31, n148_tree_31, n149_tree_31, n150_tree_31, n151_tree_31, n152_tree_31, n153_tree_31, n154_tree_31, n155_tree_31, n156_tree_31, n157_tree_31, n158_tree_31, n159_tree_31, n160_tree_31, n161_tree_31, n162_tree_31, n163_tree_31, n164_tree_31, n165_tree_31, n166_tree_31, n167_tree_31, n168_tree_31, n169_tree_31, n170_tree_31, n171_tree_31, n172_tree_31, n173_tree_31, n174_tree_31, n175_tree_31, n176_tree_31, n177_tree_31, n178_tree_31, n179_tree_31, n180_tree_31, n181_tree_31, n182_tree_31, n183_tree_31, n184_tree_31, n185_tree_31, n186_tree_31, n187_tree_31, n188_tree_31, n189_tree_31, n190_tree_31, n191_tree_31, n192_tree_31, n193_tree_31, n194_tree_31, n195_tree_31, n196_tree_31, n197_tree_31, n198_tree_31, n199_tree_31, n200_tree_31, n201_tree_31, n202_tree_31, n203_tree_31, n204_tree_31, n205_tree_31, n206_tree_31, n207_tree_31, n208_tree_31, n209_tree_31, n210_tree_31, n211_tree_31, n212_tree_31, n213_tree_31, n214_tree_31, n215_tree_31;
    assign sum[31] = n125_tree_31^n124_tree_31;
    assign n124_tree_31 = a_in[31]^b_in[31];
    assign n125_tree_31 = (n128_tree_31&n127_tree_31)|n126_tree_31;
    assign n127_tree_31 = a_in[30]|b_in[30];

    assign n126_tree_31 = a_in[30]&b_in[30];
    assign n128_tree_31 = (n131_tree_31&n130_tree_31)|n129_tree_31;
    assign n130_tree_31 = a_in[29]|b_in[29];

    assign n129_tree_31 = a_in[29]&b_in[29];
    assign n131_tree_31 = (n134_tree_31&n133_tree_31)|n132_tree_31;
    assign n133_tree_31 = a_in[28]|b_in[28];

    assign n132_tree_31 = a_in[28]&b_in[28];
    assign n134_tree_31 = (n137_tree_31&n136_tree_31)|n135_tree_31;
    assign n136_tree_31 = a_in[27]|b_in[27];

    assign n135_tree_31 = a_in[27]&b_in[27];
    assign n137_tree_31 = (n140_tree_31&n139_tree_31)|n138_tree_31;
    assign n139_tree_31 = a_in[26]|b_in[26];

    assign n138_tree_31 = a_in[26]&b_in[26];
    assign n140_tree_31 = (n143_tree_31&n142_tree_31)|n141_tree_31;
    assign n142_tree_31 = a_in[25]|b_in[25];

    assign n141_tree_31 = a_in[25]&b_in[25];
    assign n143_tree_31 = (n146_tree_31&n145_tree_31)|n144_tree_31;
    assign n145_tree_31 = a_in[24]|b_in[24];

    assign n144_tree_31 = a_in[24]&b_in[24];
    assign n146_tree_31 = (n149_tree_31&n148_tree_31)|n147_tree_31;
    assign n148_tree_31 = a_in[23]|b_in[23];

    assign n147_tree_31 = a_in[23]&b_in[23];
    assign n149_tree_31 = (n152_tree_31&n151_tree_31)|n150_tree_31;
    assign n151_tree_31 = a_in[22]|b_in[22];

    assign n150_tree_31 = a_in[22]&b_in[22];
    assign n152_tree_31 = (n155_tree_31&n154_tree_31)|n153_tree_31;
    assign n154_tree_31 = a_in[21]|b_in[21];

    assign n153_tree_31 = a_in[21]&b_in[21];
    assign n155_tree_31 = (n158_tree_31&n157_tree_31)|n156_tree_31;
    assign n157_tree_31 = a_in[20]|b_in[20];

    assign n156_tree_31 = a_in[20]&b_in[20];
    assign n158_tree_31 = (n161_tree_31&n160_tree_31)|n159_tree_31;
    assign n160_tree_31 = a_in[19]|b_in[19];

    assign n159_tree_31 = a_in[19]&b_in[19];
    assign n161_tree_31 = (n164_tree_31&n163_tree_31)|n162_tree_31;
    assign n163_tree_31 = a_in[18]|b_in[18];

    assign n162_tree_31 = a_in[18]&b_in[18];
    assign n164_tree_31 = (n167_tree_31&n166_tree_31)|n165_tree_31;
    assign n166_tree_31 = a_in[17]|b_in[17];

    assign n165_tree_31 = a_in[17]&b_in[17];
    assign n167_tree_31 = (n170_tree_31&n169_tree_31)|n168_tree_31;
    assign n169_tree_31 = a_in[16]|b_in[16];

    assign n168_tree_31 = a_in[16]&b_in[16];
    assign n170_tree_31 = (n173_tree_31&n172_tree_31)|n171_tree_31;
    assign n172_tree_31 = a_in[15]|b_in[15];

    assign n171_tree_31 = a_in[15]&b_in[15];
    assign n173_tree_31 = (n176_tree_31&n175_tree_31)|n174_tree_31;
    assign n175_tree_31 = a_in[14]|b_in[14];

    assign n174_tree_31 = a_in[14]&b_in[14];
    assign n176_tree_31 = (n179_tree_31&n178_tree_31)|n177_tree_31;
    assign n178_tree_31 = a_in[13]|b_in[13];

    assign n177_tree_31 = a_in[13]&b_in[13];
    assign n179_tree_31 = (n182_tree_31&n181_tree_31)|n180_tree_31;
    assign n181_tree_31 = a_in[12]|b_in[12];

    assign n180_tree_31 = a_in[12]&b_in[12];
    assign n182_tree_31 = (n185_tree_31&n184_tree_31)|n183_tree_31;
    assign n184_tree_31 = a_in[11]|b_in[11];

    assign n183_tree_31 = a_in[11]&b_in[11];
    assign n185_tree_31 = (n188_tree_31&n187_tree_31)|n186_tree_31;
    assign n187_tree_31 = a_in[10]|b_in[10];

    assign n186_tree_31 = a_in[10]&b_in[10];
    assign n188_tree_31 = (n191_tree_31&n190_tree_31)|n189_tree_31;
    assign n190_tree_31 = a_in[9]|b_in[9];

    assign n189_tree_31 = a_in[9]&b_in[9];
    assign n191_tree_31 = (n194_tree_31&n193_tree_31)|n192_tree_31;
    assign n193_tree_31 = a_in[8]|b_in[8];

    assign n192_tree_31 = a_in[8]&b_in[8];
    assign n194_tree_31 = (n197_tree_31&n196_tree_31)|n195_tree_31;
    assign n196_tree_31 = a_in[7]|b_in[7];

    assign n195_tree_31 = a_in[7]&b_in[7];
    assign n197_tree_31 = (n200_tree_31&n199_tree_31)|n198_tree_31;
    assign n199_tree_31 = a_in[6]|b_in[6];

    assign n198_tree_31 = a_in[6]&b_in[6];
    assign n200_tree_31 = (n203_tree_31&n202_tree_31)|n201_tree_31;
    assign n202_tree_31 = a_in[5]|b_in[5];

    assign n201_tree_31 = a_in[5]&b_in[5];
    assign n203_tree_31 = (n206_tree_31&n205_tree_31)|n204_tree_31;
    assign n205_tree_31 = a_in[4]|b_in[4];

    assign n204_tree_31 = a_in[4]&b_in[4];
    assign n206_tree_31 = (n209_tree_31&n208_tree_31)|n207_tree_31;
    assign n208_tree_31 = a_in[3]|b_in[3];

    assign n207_tree_31 = a_in[3]&b_in[3];
    assign n209_tree_31 = (n212_tree_31&n211_tree_31)|n210_tree_31;
    assign n211_tree_31 = a_in[2]|b_in[2];

    assign n210_tree_31 = a_in[2]&b_in[2];
    assign n212_tree_31 = (n215_tree_31&n214_tree_31)|n213_tree_31;
    assign n214_tree_31 = a_in[1]|b_in[1];

    assign n213_tree_31 = a_in[1]&b_in[1];
    assign n215_tree_31 = a_in[0]&b_in[0];

// adder_forest tree_30
	wire n120_tree_30, n121_tree_30, n122_tree_30, n123_tree_30, n124_tree_30, n125_tree_30, n126_tree_30, n127_tree_30, n128_tree_30, n129_tree_30, n130_tree_30, n131_tree_30, n132_tree_30, n133_tree_30, n134_tree_30, n135_tree_30, n136_tree_30, n137_tree_30, n138_tree_30, n139_tree_30, n140_tree_30, n141_tree_30, n142_tree_30, n143_tree_30, n144_tree_30, n145_tree_30, n146_tree_30, n147_tree_30, n148_tree_30, n149_tree_30, n150_tree_30, n151_tree_30, n152_tree_30, n153_tree_30, n154_tree_30, n155_tree_30, n156_tree_30, n157_tree_30, n158_tree_30, n159_tree_30, n160_tree_30, n161_tree_30, n162_tree_30, n163_tree_30, n164_tree_30, n165_tree_30, n166_tree_30, n167_tree_30, n168_tree_30, n169_tree_30, n170_tree_30, n171_tree_30, n172_tree_30, n173_tree_30, n174_tree_30, n175_tree_30, n176_tree_30, n177_tree_30, n178_tree_30, n179_tree_30, n180_tree_30, n181_tree_30, n182_tree_30, n183_tree_30, n184_tree_30, n185_tree_30, n186_tree_30, n187_tree_30, n188_tree_30, n189_tree_30, n190_tree_30, n191_tree_30, n192_tree_30, n193_tree_30, n194_tree_30, n195_tree_30, n196_tree_30, n197_tree_30, n198_tree_30, n199_tree_30, n200_tree_30, n201_tree_30, n202_tree_30, n203_tree_30, n204_tree_30, n205_tree_30, n206_tree_30, n207_tree_30, n208_tree_30;
    assign sum[30] = n121_tree_30^n120_tree_30;
    assign n120_tree_30 = a_in[30]^b_in[30];
    assign n121_tree_30 = (n124_tree_30&n123_tree_30)|n122_tree_30;
    assign n123_tree_30 = a_in[29]|b_in[29];

    assign n122_tree_30 = a_in[29]&b_in[29];
    assign n124_tree_30 = (n127_tree_30&n126_tree_30)|n125_tree_30;
    assign n126_tree_30 = a_in[28]|b_in[28];

    assign n125_tree_30 = a_in[28]&b_in[28];
    assign n127_tree_30 = (n130_tree_30&n129_tree_30)|n128_tree_30;
    assign n129_tree_30 = a_in[27]|b_in[27];

    assign n128_tree_30 = a_in[27]&b_in[27];
    assign n130_tree_30 = (n133_tree_30&n132_tree_30)|n131_tree_30;
    assign n132_tree_30 = a_in[26]|b_in[26];

    assign n131_tree_30 = a_in[26]&b_in[26];
    assign n133_tree_30 = (n136_tree_30&n135_tree_30)|n134_tree_30;
    assign n135_tree_30 = a_in[25]|b_in[25];

    assign n134_tree_30 = a_in[25]&b_in[25];
    assign n136_tree_30 = (n139_tree_30&n138_tree_30)|n137_tree_30;
    assign n138_tree_30 = a_in[24]|b_in[24];

    assign n137_tree_30 = a_in[24]&b_in[24];
    assign n139_tree_30 = (n142_tree_30&n141_tree_30)|n140_tree_30;
    assign n141_tree_30 = a_in[23]|b_in[23];

    assign n140_tree_30 = a_in[23]&b_in[23];
    assign n142_tree_30 = (n145_tree_30&n144_tree_30)|n143_tree_30;
    assign n144_tree_30 = a_in[22]|b_in[22];

    assign n143_tree_30 = a_in[22]&b_in[22];
    assign n145_tree_30 = (n148_tree_30&n147_tree_30)|n146_tree_30;
    assign n147_tree_30 = a_in[21]|b_in[21];

    assign n146_tree_30 = a_in[21]&b_in[21];
    assign n148_tree_30 = (n151_tree_30&n150_tree_30)|n149_tree_30;
    assign n150_tree_30 = a_in[20]|b_in[20];

    assign n149_tree_30 = a_in[20]&b_in[20];
    assign n151_tree_30 = (n154_tree_30&n153_tree_30)|n152_tree_30;
    assign n153_tree_30 = a_in[19]|b_in[19];

    assign n152_tree_30 = a_in[19]&b_in[19];
    assign n154_tree_30 = (n157_tree_30&n156_tree_30)|n155_tree_30;
    assign n156_tree_30 = a_in[18]|b_in[18];

    assign n155_tree_30 = a_in[18]&b_in[18];
    assign n157_tree_30 = (n160_tree_30&n159_tree_30)|n158_tree_30;
    assign n159_tree_30 = a_in[17]|b_in[17];

    assign n158_tree_30 = a_in[17]&b_in[17];
    assign n160_tree_30 = (n163_tree_30&n162_tree_30)|n161_tree_30;
    assign n162_tree_30 = a_in[16]|b_in[16];

    assign n161_tree_30 = a_in[16]&b_in[16];
    assign n163_tree_30 = (n166_tree_30&n165_tree_30)|n164_tree_30;
    assign n165_tree_30 = a_in[15]|b_in[15];

    assign n164_tree_30 = a_in[15]&b_in[15];
    assign n166_tree_30 = (n169_tree_30&n168_tree_30)|n167_tree_30;
    assign n168_tree_30 = a_in[14]|b_in[14];

    assign n167_tree_30 = a_in[14]&b_in[14];
    assign n169_tree_30 = (n172_tree_30&n171_tree_30)|n170_tree_30;
    assign n171_tree_30 = a_in[13]|b_in[13];

    assign n170_tree_30 = a_in[13]&b_in[13];
    assign n172_tree_30 = (n175_tree_30&n174_tree_30)|n173_tree_30;
    assign n174_tree_30 = a_in[12]|b_in[12];

    assign n173_tree_30 = a_in[12]&b_in[12];
    assign n175_tree_30 = (n178_tree_30&n177_tree_30)|n176_tree_30;
    assign n177_tree_30 = a_in[11]|b_in[11];

    assign n176_tree_30 = a_in[11]&b_in[11];
    assign n178_tree_30 = (n181_tree_30&n180_tree_30)|n179_tree_30;
    assign n180_tree_30 = a_in[10]|b_in[10];

    assign n179_tree_30 = a_in[10]&b_in[10];
    assign n181_tree_30 = (n184_tree_30&n183_tree_30)|n182_tree_30;
    assign n183_tree_30 = a_in[9]|b_in[9];

    assign n182_tree_30 = a_in[9]&b_in[9];
    assign n184_tree_30 = (n187_tree_30&n186_tree_30)|n185_tree_30;
    assign n186_tree_30 = a_in[8]|b_in[8];

    assign n185_tree_30 = a_in[8]&b_in[8];
    assign n187_tree_30 = (n190_tree_30&n189_tree_30)|n188_tree_30;
    assign n189_tree_30 = a_in[7]|b_in[7];

    assign n188_tree_30 = a_in[7]&b_in[7];
    assign n190_tree_30 = (n193_tree_30&n192_tree_30)|n191_tree_30;
    assign n192_tree_30 = a_in[6]|b_in[6];

    assign n191_tree_30 = a_in[6]&b_in[6];
    assign n193_tree_30 = (n196_tree_30&n195_tree_30)|n194_tree_30;
    assign n195_tree_30 = a_in[5]|b_in[5];

    assign n194_tree_30 = a_in[5]&b_in[5];
    assign n196_tree_30 = (n199_tree_30&n198_tree_30)|n197_tree_30;
    assign n198_tree_30 = a_in[4]|b_in[4];

    assign n197_tree_30 = a_in[4]&b_in[4];
    assign n199_tree_30 = (n202_tree_30&n201_tree_30)|n200_tree_30;
    assign n201_tree_30 = a_in[3]|b_in[3];

    assign n200_tree_30 = a_in[3]&b_in[3];
    assign n202_tree_30 = (n205_tree_30&n204_tree_30)|n203_tree_30;
    assign n204_tree_30 = a_in[2]|b_in[2];

    assign n203_tree_30 = a_in[2]&b_in[2];
    assign n205_tree_30 = (n208_tree_30&n207_tree_30)|n206_tree_30;
    assign n207_tree_30 = a_in[1]|b_in[1];

    assign n206_tree_30 = a_in[1]&b_in[1];
    assign n208_tree_30 = a_in[0]&b_in[0];

// adder_forest tree_29
	wire n116_tree_29, n117_tree_29, n118_tree_29, n119_tree_29, n120_tree_29, n121_tree_29, n122_tree_29, n123_tree_29, n124_tree_29, n125_tree_29, n126_tree_29, n127_tree_29, n128_tree_29, n129_tree_29, n130_tree_29, n131_tree_29, n132_tree_29, n133_tree_29, n134_tree_29, n135_tree_29, n136_tree_29, n137_tree_29, n138_tree_29, n139_tree_29, n140_tree_29, n141_tree_29, n142_tree_29, n143_tree_29, n144_tree_29, n145_tree_29, n146_tree_29, n147_tree_29, n148_tree_29, n149_tree_29, n150_tree_29, n151_tree_29, n152_tree_29, n153_tree_29, n154_tree_29, n155_tree_29, n156_tree_29, n157_tree_29, n158_tree_29, n159_tree_29, n160_tree_29, n161_tree_29, n162_tree_29, n163_tree_29, n164_tree_29, n165_tree_29, n166_tree_29, n167_tree_29, n168_tree_29, n169_tree_29, n170_tree_29, n171_tree_29, n172_tree_29, n173_tree_29, n174_tree_29, n175_tree_29, n176_tree_29, n177_tree_29, n178_tree_29, n179_tree_29, n180_tree_29, n181_tree_29, n182_tree_29, n183_tree_29, n184_tree_29, n185_tree_29, n186_tree_29, n187_tree_29, n188_tree_29, n189_tree_29, n190_tree_29, n191_tree_29, n192_tree_29, n193_tree_29, n194_tree_29, n195_tree_29, n196_tree_29, n197_tree_29, n198_tree_29, n199_tree_29, n200_tree_29, n201_tree_29;
    assign sum[29] = n117_tree_29^n116_tree_29;
    assign n116_tree_29 = a_in[29]^b_in[29];
    assign n117_tree_29 = (n120_tree_29&n119_tree_29)|n118_tree_29;
    assign n119_tree_29 = a_in[28]|b_in[28];

    assign n118_tree_29 = a_in[28]&b_in[28];
    assign n120_tree_29 = (n123_tree_29&n122_tree_29)|n121_tree_29;
    assign n122_tree_29 = a_in[27]|b_in[27];

    assign n121_tree_29 = a_in[27]&b_in[27];
    assign n123_tree_29 = (n126_tree_29&n125_tree_29)|n124_tree_29;
    assign n125_tree_29 = a_in[26]|b_in[26];

    assign n124_tree_29 = a_in[26]&b_in[26];
    assign n126_tree_29 = (n129_tree_29&n128_tree_29)|n127_tree_29;
    assign n128_tree_29 = a_in[25]|b_in[25];

    assign n127_tree_29 = a_in[25]&b_in[25];
    assign n129_tree_29 = (n132_tree_29&n131_tree_29)|n130_tree_29;
    assign n131_tree_29 = a_in[24]|b_in[24];

    assign n130_tree_29 = a_in[24]&b_in[24];
    assign n132_tree_29 = (n135_tree_29&n134_tree_29)|n133_tree_29;
    assign n134_tree_29 = a_in[23]|b_in[23];

    assign n133_tree_29 = a_in[23]&b_in[23];
    assign n135_tree_29 = (n138_tree_29&n137_tree_29)|n136_tree_29;
    assign n137_tree_29 = a_in[22]|b_in[22];

    assign n136_tree_29 = a_in[22]&b_in[22];
    assign n138_tree_29 = (n141_tree_29&n140_tree_29)|n139_tree_29;
    assign n140_tree_29 = a_in[21]|b_in[21];

    assign n139_tree_29 = a_in[21]&b_in[21];
    assign n141_tree_29 = (n144_tree_29&n143_tree_29)|n142_tree_29;
    assign n143_tree_29 = a_in[20]|b_in[20];

    assign n142_tree_29 = a_in[20]&b_in[20];
    assign n144_tree_29 = (n147_tree_29&n146_tree_29)|n145_tree_29;
    assign n146_tree_29 = a_in[19]|b_in[19];

    assign n145_tree_29 = a_in[19]&b_in[19];
    assign n147_tree_29 = (n150_tree_29&n149_tree_29)|n148_tree_29;
    assign n149_tree_29 = a_in[18]|b_in[18];

    assign n148_tree_29 = a_in[18]&b_in[18];
    assign n150_tree_29 = (n153_tree_29&n152_tree_29)|n151_tree_29;
    assign n152_tree_29 = a_in[17]|b_in[17];

    assign n151_tree_29 = a_in[17]&b_in[17];
    assign n153_tree_29 = (n156_tree_29&n155_tree_29)|n154_tree_29;
    assign n155_tree_29 = a_in[16]|b_in[16];

    assign n154_tree_29 = a_in[16]&b_in[16];
    assign n156_tree_29 = (n159_tree_29&n158_tree_29)|n157_tree_29;
    assign n158_tree_29 = a_in[15]|b_in[15];

    assign n157_tree_29 = a_in[15]&b_in[15];
    assign n159_tree_29 = (n162_tree_29&n161_tree_29)|n160_tree_29;
    assign n161_tree_29 = a_in[14]|b_in[14];

    assign n160_tree_29 = a_in[14]&b_in[14];
    assign n162_tree_29 = (n165_tree_29&n164_tree_29)|n163_tree_29;
    assign n164_tree_29 = a_in[13]|b_in[13];

    assign n163_tree_29 = a_in[13]&b_in[13];
    assign n165_tree_29 = (n168_tree_29&n167_tree_29)|n166_tree_29;
    assign n167_tree_29 = a_in[12]|b_in[12];

    assign n166_tree_29 = a_in[12]&b_in[12];
    assign n168_tree_29 = (n171_tree_29&n170_tree_29)|n169_tree_29;
    assign n170_tree_29 = a_in[11]|b_in[11];

    assign n169_tree_29 = a_in[11]&b_in[11];
    assign n171_tree_29 = (n174_tree_29&n173_tree_29)|n172_tree_29;
    assign n173_tree_29 = a_in[10]|b_in[10];

    assign n172_tree_29 = a_in[10]&b_in[10];
    assign n174_tree_29 = (n177_tree_29&n176_tree_29)|n175_tree_29;
    assign n176_tree_29 = a_in[9]|b_in[9];

    assign n175_tree_29 = a_in[9]&b_in[9];
    assign n177_tree_29 = (n180_tree_29&n179_tree_29)|n178_tree_29;
    assign n179_tree_29 = a_in[8]|b_in[8];

    assign n178_tree_29 = a_in[8]&b_in[8];
    assign n180_tree_29 = (n183_tree_29&n182_tree_29)|n181_tree_29;
    assign n182_tree_29 = a_in[7]|b_in[7];

    assign n181_tree_29 = a_in[7]&b_in[7];
    assign n183_tree_29 = (n186_tree_29&n185_tree_29)|n184_tree_29;
    assign n185_tree_29 = a_in[6]|b_in[6];

    assign n184_tree_29 = a_in[6]&b_in[6];
    assign n186_tree_29 = (n189_tree_29&n188_tree_29)|n187_tree_29;
    assign n188_tree_29 = a_in[5]|b_in[5];

    assign n187_tree_29 = a_in[5]&b_in[5];
    assign n189_tree_29 = (n192_tree_29&n191_tree_29)|n190_tree_29;
    assign n191_tree_29 = a_in[4]|b_in[4];

    assign n190_tree_29 = a_in[4]&b_in[4];
    assign n192_tree_29 = (n195_tree_29&n194_tree_29)|n193_tree_29;
    assign n194_tree_29 = a_in[3]|b_in[3];

    assign n193_tree_29 = a_in[3]&b_in[3];
    assign n195_tree_29 = (n198_tree_29&n197_tree_29)|n196_tree_29;
    assign n197_tree_29 = a_in[2]|b_in[2];

    assign n196_tree_29 = a_in[2]&b_in[2];
    assign n198_tree_29 = (n201_tree_29&n200_tree_29)|n199_tree_29;
    assign n200_tree_29 = a_in[1]|b_in[1];

    assign n199_tree_29 = a_in[1]&b_in[1];
    assign n201_tree_29 = a_in[0]&b_in[0];

// adder_forest tree_28
	wire n112_tree_28, n113_tree_28, n114_tree_28, n115_tree_28, n116_tree_28, n117_tree_28, n118_tree_28, n119_tree_28, n120_tree_28, n121_tree_28, n122_tree_28, n123_tree_28, n124_tree_28, n125_tree_28, n126_tree_28, n127_tree_28, n128_tree_28, n129_tree_28, n130_tree_28, n131_tree_28, n132_tree_28, n133_tree_28, n134_tree_28, n135_tree_28, n136_tree_28, n137_tree_28, n138_tree_28, n139_tree_28, n140_tree_28, n141_tree_28, n142_tree_28, n143_tree_28, n144_tree_28, n145_tree_28, n146_tree_28, n147_tree_28, n148_tree_28, n149_tree_28, n150_tree_28, n151_tree_28, n152_tree_28, n153_tree_28, n154_tree_28, n155_tree_28, n156_tree_28, n157_tree_28, n158_tree_28, n159_tree_28, n160_tree_28, n161_tree_28, n162_tree_28, n163_tree_28, n164_tree_28, n165_tree_28, n166_tree_28, n167_tree_28, n168_tree_28, n169_tree_28, n170_tree_28, n171_tree_28, n172_tree_28, n173_tree_28, n174_tree_28, n175_tree_28, n176_tree_28, n177_tree_28, n178_tree_28, n179_tree_28, n180_tree_28, n181_tree_28, n182_tree_28, n183_tree_28, n184_tree_28, n185_tree_28, n186_tree_28, n187_tree_28, n188_tree_28, n189_tree_28, n190_tree_28, n191_tree_28, n192_tree_28, n193_tree_28, n194_tree_28;
    assign sum[28] = n113_tree_28^n112_tree_28;
    assign n112_tree_28 = a_in[28]^b_in[28];
    assign n113_tree_28 = (n116_tree_28&n115_tree_28)|n114_tree_28;
    assign n115_tree_28 = a_in[27]|b_in[27];

    assign n114_tree_28 = a_in[27]&b_in[27];
    assign n116_tree_28 = (n119_tree_28&n118_tree_28)|n117_tree_28;
    assign n118_tree_28 = a_in[26]|b_in[26];

    assign n117_tree_28 = a_in[26]&b_in[26];
    assign n119_tree_28 = (n122_tree_28&n121_tree_28)|n120_tree_28;
    assign n121_tree_28 = a_in[25]|b_in[25];

    assign n120_tree_28 = a_in[25]&b_in[25];
    assign n122_tree_28 = (n125_tree_28&n124_tree_28)|n123_tree_28;
    assign n124_tree_28 = a_in[24]|b_in[24];

    assign n123_tree_28 = a_in[24]&b_in[24];
    assign n125_tree_28 = (n128_tree_28&n127_tree_28)|n126_tree_28;
    assign n127_tree_28 = a_in[23]|b_in[23];

    assign n126_tree_28 = a_in[23]&b_in[23];
    assign n128_tree_28 = (n131_tree_28&n130_tree_28)|n129_tree_28;
    assign n130_tree_28 = a_in[22]|b_in[22];

    assign n129_tree_28 = a_in[22]&b_in[22];
    assign n131_tree_28 = (n134_tree_28&n133_tree_28)|n132_tree_28;
    assign n133_tree_28 = a_in[21]|b_in[21];

    assign n132_tree_28 = a_in[21]&b_in[21];
    assign n134_tree_28 = (n137_tree_28&n136_tree_28)|n135_tree_28;
    assign n136_tree_28 = a_in[20]|b_in[20];

    assign n135_tree_28 = a_in[20]&b_in[20];
    assign n137_tree_28 = (n140_tree_28&n139_tree_28)|n138_tree_28;
    assign n139_tree_28 = a_in[19]|b_in[19];

    assign n138_tree_28 = a_in[19]&b_in[19];
    assign n140_tree_28 = (n143_tree_28&n142_tree_28)|n141_tree_28;
    assign n142_tree_28 = a_in[18]|b_in[18];

    assign n141_tree_28 = a_in[18]&b_in[18];
    assign n143_tree_28 = (n146_tree_28&n145_tree_28)|n144_tree_28;
    assign n145_tree_28 = a_in[17]|b_in[17];

    assign n144_tree_28 = a_in[17]&b_in[17];
    assign n146_tree_28 = (n149_tree_28&n148_tree_28)|n147_tree_28;
    assign n148_tree_28 = a_in[16]|b_in[16];

    assign n147_tree_28 = a_in[16]&b_in[16];
    assign n149_tree_28 = (n152_tree_28&n151_tree_28)|n150_tree_28;
    assign n151_tree_28 = a_in[15]|b_in[15];

    assign n150_tree_28 = a_in[15]&b_in[15];
    assign n152_tree_28 = (n155_tree_28&n154_tree_28)|n153_tree_28;
    assign n154_tree_28 = a_in[14]|b_in[14];

    assign n153_tree_28 = a_in[14]&b_in[14];
    assign n155_tree_28 = (n158_tree_28&n157_tree_28)|n156_tree_28;
    assign n157_tree_28 = a_in[13]|b_in[13];

    assign n156_tree_28 = a_in[13]&b_in[13];
    assign n158_tree_28 = (n161_tree_28&n160_tree_28)|n159_tree_28;
    assign n160_tree_28 = a_in[12]|b_in[12];

    assign n159_tree_28 = a_in[12]&b_in[12];
    assign n161_tree_28 = (n164_tree_28&n163_tree_28)|n162_tree_28;
    assign n163_tree_28 = a_in[11]|b_in[11];

    assign n162_tree_28 = a_in[11]&b_in[11];
    assign n164_tree_28 = (n167_tree_28&n166_tree_28)|n165_tree_28;
    assign n166_tree_28 = a_in[10]|b_in[10];

    assign n165_tree_28 = a_in[10]&b_in[10];
    assign n167_tree_28 = (n170_tree_28&n169_tree_28)|n168_tree_28;
    assign n169_tree_28 = a_in[9]|b_in[9];

    assign n168_tree_28 = a_in[9]&b_in[9];
    assign n170_tree_28 = (n173_tree_28&n172_tree_28)|n171_tree_28;
    assign n172_tree_28 = a_in[8]|b_in[8];

    assign n171_tree_28 = a_in[8]&b_in[8];
    assign n173_tree_28 = (n176_tree_28&n175_tree_28)|n174_tree_28;
    assign n175_tree_28 = a_in[7]|b_in[7];

    assign n174_tree_28 = a_in[7]&b_in[7];
    assign n176_tree_28 = (n179_tree_28&n178_tree_28)|n177_tree_28;
    assign n178_tree_28 = a_in[6]|b_in[6];

    assign n177_tree_28 = a_in[6]&b_in[6];
    assign n179_tree_28 = (n182_tree_28&n181_tree_28)|n180_tree_28;
    assign n181_tree_28 = a_in[5]|b_in[5];

    assign n180_tree_28 = a_in[5]&b_in[5];
    assign n182_tree_28 = (n185_tree_28&n184_tree_28)|n183_tree_28;
    assign n184_tree_28 = a_in[4]|b_in[4];

    assign n183_tree_28 = a_in[4]&b_in[4];
    assign n185_tree_28 = (n188_tree_28&n187_tree_28)|n186_tree_28;
    assign n187_tree_28 = a_in[3]|b_in[3];

    assign n186_tree_28 = a_in[3]&b_in[3];
    assign n188_tree_28 = (n191_tree_28&n190_tree_28)|n189_tree_28;
    assign n190_tree_28 = a_in[2]|b_in[2];

    assign n189_tree_28 = a_in[2]&b_in[2];
    assign n191_tree_28 = (n194_tree_28&n193_tree_28)|n192_tree_28;
    assign n193_tree_28 = a_in[1]|b_in[1];

    assign n192_tree_28 = a_in[1]&b_in[1];
    assign n194_tree_28 = a_in[0]&b_in[0];

// adder_forest tree_27
	wire n108_tree_27, n109_tree_27, n110_tree_27, n111_tree_27, n112_tree_27, n113_tree_27, n114_tree_27, n115_tree_27, n116_tree_27, n117_tree_27, n118_tree_27, n119_tree_27, n120_tree_27, n121_tree_27, n122_tree_27, n123_tree_27, n124_tree_27, n125_tree_27, n126_tree_27, n127_tree_27, n128_tree_27, n129_tree_27, n130_tree_27, n131_tree_27, n132_tree_27, n133_tree_27, n134_tree_27, n135_tree_27, n136_tree_27, n137_tree_27, n138_tree_27, n139_tree_27, n140_tree_27, n141_tree_27, n142_tree_27, n143_tree_27, n144_tree_27, n145_tree_27, n146_tree_27, n147_tree_27, n148_tree_27, n149_tree_27, n150_tree_27, n151_tree_27, n152_tree_27, n153_tree_27, n154_tree_27, n155_tree_27, n156_tree_27, n157_tree_27, n158_tree_27, n159_tree_27, n160_tree_27, n161_tree_27, n162_tree_27, n163_tree_27, n164_tree_27, n165_tree_27, n166_tree_27, n167_tree_27, n168_tree_27, n169_tree_27, n170_tree_27, n171_tree_27, n172_tree_27, n173_tree_27, n174_tree_27, n175_tree_27, n176_tree_27, n177_tree_27, n178_tree_27, n179_tree_27, n180_tree_27, n181_tree_27, n182_tree_27, n183_tree_27, n184_tree_27, n185_tree_27, n186_tree_27, n187_tree_27;
    assign sum[27] = n109_tree_27^n108_tree_27;
    assign n108_tree_27 = a_in[27]^b_in[27];
    assign n109_tree_27 = (n112_tree_27&n111_tree_27)|n110_tree_27;
    assign n111_tree_27 = a_in[26]|b_in[26];

    assign n110_tree_27 = a_in[26]&b_in[26];
    assign n112_tree_27 = (n115_tree_27&n114_tree_27)|n113_tree_27;
    assign n114_tree_27 = a_in[25]|b_in[25];

    assign n113_tree_27 = a_in[25]&b_in[25];
    assign n115_tree_27 = (n118_tree_27&n117_tree_27)|n116_tree_27;
    assign n117_tree_27 = a_in[24]|b_in[24];

    assign n116_tree_27 = a_in[24]&b_in[24];
    assign n118_tree_27 = (n121_tree_27&n120_tree_27)|n119_tree_27;
    assign n120_tree_27 = a_in[23]|b_in[23];

    assign n119_tree_27 = a_in[23]&b_in[23];
    assign n121_tree_27 = (n124_tree_27&n123_tree_27)|n122_tree_27;
    assign n123_tree_27 = a_in[22]|b_in[22];

    assign n122_tree_27 = a_in[22]&b_in[22];
    assign n124_tree_27 = (n127_tree_27&n126_tree_27)|n125_tree_27;
    assign n126_tree_27 = a_in[21]|b_in[21];

    assign n125_tree_27 = a_in[21]&b_in[21];
    assign n127_tree_27 = (n130_tree_27&n129_tree_27)|n128_tree_27;
    assign n129_tree_27 = a_in[20]|b_in[20];

    assign n128_tree_27 = a_in[20]&b_in[20];
    assign n130_tree_27 = (n133_tree_27&n132_tree_27)|n131_tree_27;
    assign n132_tree_27 = a_in[19]|b_in[19];

    assign n131_tree_27 = a_in[19]&b_in[19];
    assign n133_tree_27 = (n136_tree_27&n135_tree_27)|n134_tree_27;
    assign n135_tree_27 = a_in[18]|b_in[18];

    assign n134_tree_27 = a_in[18]&b_in[18];
    assign n136_tree_27 = (n139_tree_27&n138_tree_27)|n137_tree_27;
    assign n138_tree_27 = a_in[17]|b_in[17];

    assign n137_tree_27 = a_in[17]&b_in[17];
    assign n139_tree_27 = (n142_tree_27&n141_tree_27)|n140_tree_27;
    assign n141_tree_27 = a_in[16]|b_in[16];

    assign n140_tree_27 = a_in[16]&b_in[16];
    assign n142_tree_27 = (n145_tree_27&n144_tree_27)|n143_tree_27;
    assign n144_tree_27 = a_in[15]|b_in[15];

    assign n143_tree_27 = a_in[15]&b_in[15];
    assign n145_tree_27 = (n148_tree_27&n147_tree_27)|n146_tree_27;
    assign n147_tree_27 = a_in[14]|b_in[14];

    assign n146_tree_27 = a_in[14]&b_in[14];
    assign n148_tree_27 = (n151_tree_27&n150_tree_27)|n149_tree_27;
    assign n150_tree_27 = a_in[13]|b_in[13];

    assign n149_tree_27 = a_in[13]&b_in[13];
    assign n151_tree_27 = (n154_tree_27&n153_tree_27)|n152_tree_27;
    assign n153_tree_27 = a_in[12]|b_in[12];

    assign n152_tree_27 = a_in[12]&b_in[12];
    assign n154_tree_27 = (n157_tree_27&n156_tree_27)|n155_tree_27;
    assign n156_tree_27 = a_in[11]|b_in[11];

    assign n155_tree_27 = a_in[11]&b_in[11];
    assign n157_tree_27 = (n160_tree_27&n159_tree_27)|n158_tree_27;
    assign n159_tree_27 = a_in[10]|b_in[10];

    assign n158_tree_27 = a_in[10]&b_in[10];
    assign n160_tree_27 = (n163_tree_27&n162_tree_27)|n161_tree_27;
    assign n162_tree_27 = a_in[9]|b_in[9];

    assign n161_tree_27 = a_in[9]&b_in[9];
    assign n163_tree_27 = (n166_tree_27&n165_tree_27)|n164_tree_27;
    assign n165_tree_27 = a_in[8]|b_in[8];

    assign n164_tree_27 = a_in[8]&b_in[8];
    assign n166_tree_27 = (n169_tree_27&n168_tree_27)|n167_tree_27;
    assign n168_tree_27 = a_in[7]|b_in[7];

    assign n167_tree_27 = a_in[7]&b_in[7];
    assign n169_tree_27 = (n172_tree_27&n171_tree_27)|n170_tree_27;
    assign n171_tree_27 = a_in[6]|b_in[6];

    assign n170_tree_27 = a_in[6]&b_in[6];
    assign n172_tree_27 = (n175_tree_27&n174_tree_27)|n173_tree_27;
    assign n174_tree_27 = a_in[5]|b_in[5];

    assign n173_tree_27 = a_in[5]&b_in[5];
    assign n175_tree_27 = (n178_tree_27&n177_tree_27)|n176_tree_27;
    assign n177_tree_27 = a_in[4]|b_in[4];

    assign n176_tree_27 = a_in[4]&b_in[4];
    assign n178_tree_27 = (n181_tree_27&n180_tree_27)|n179_tree_27;
    assign n180_tree_27 = a_in[3]|b_in[3];

    assign n179_tree_27 = a_in[3]&b_in[3];
    assign n181_tree_27 = (n184_tree_27&n183_tree_27)|n182_tree_27;
    assign n183_tree_27 = a_in[2]|b_in[2];

    assign n182_tree_27 = a_in[2]&b_in[2];
    assign n184_tree_27 = (n187_tree_27&n186_tree_27)|n185_tree_27;
    assign n186_tree_27 = a_in[1]|b_in[1];

    assign n185_tree_27 = a_in[1]&b_in[1];
    assign n187_tree_27 = a_in[0]&b_in[0];

// adder_forest tree_26
	wire n104_tree_26, n105_tree_26, n106_tree_26, n107_tree_26, n108_tree_26, n109_tree_26, n110_tree_26, n111_tree_26, n112_tree_26, n113_tree_26, n114_tree_26, n115_tree_26, n116_tree_26, n117_tree_26, n118_tree_26, n119_tree_26, n120_tree_26, n121_tree_26, n122_tree_26, n123_tree_26, n124_tree_26, n125_tree_26, n126_tree_26, n127_tree_26, n128_tree_26, n129_tree_26, n130_tree_26, n131_tree_26, n132_tree_26, n133_tree_26, n134_tree_26, n135_tree_26, n136_tree_26, n137_tree_26, n138_tree_26, n139_tree_26, n140_tree_26, n141_tree_26, n142_tree_26, n143_tree_26, n144_tree_26, n145_tree_26, n146_tree_26, n147_tree_26, n148_tree_26, n149_tree_26, n150_tree_26, n151_tree_26, n152_tree_26, n153_tree_26, n154_tree_26, n155_tree_26, n156_tree_26, n157_tree_26, n158_tree_26, n159_tree_26, n160_tree_26, n161_tree_26, n162_tree_26, n163_tree_26, n164_tree_26, n165_tree_26, n166_tree_26, n167_tree_26, n168_tree_26, n169_tree_26, n170_tree_26, n171_tree_26, n172_tree_26, n173_tree_26, n174_tree_26, n175_tree_26, n176_tree_26, n177_tree_26, n178_tree_26, n179_tree_26, n180_tree_26;
    assign sum[26] = n105_tree_26^n104_tree_26;
    assign n104_tree_26 = a_in[26]^b_in[26];
    assign n105_tree_26 = (n108_tree_26&n107_tree_26)|n106_tree_26;
    assign n107_tree_26 = a_in[25]|b_in[25];

    assign n106_tree_26 = a_in[25]&b_in[25];
    assign n108_tree_26 = (n111_tree_26&n110_tree_26)|n109_tree_26;
    assign n110_tree_26 = a_in[24]|b_in[24];

    assign n109_tree_26 = a_in[24]&b_in[24];
    assign n111_tree_26 = (n114_tree_26&n113_tree_26)|n112_tree_26;
    assign n113_tree_26 = a_in[23]|b_in[23];

    assign n112_tree_26 = a_in[23]&b_in[23];
    assign n114_tree_26 = (n117_tree_26&n116_tree_26)|n115_tree_26;
    assign n116_tree_26 = a_in[22]|b_in[22];

    assign n115_tree_26 = a_in[22]&b_in[22];
    assign n117_tree_26 = (n120_tree_26&n119_tree_26)|n118_tree_26;
    assign n119_tree_26 = a_in[21]|b_in[21];

    assign n118_tree_26 = a_in[21]&b_in[21];
    assign n120_tree_26 = (n123_tree_26&n122_tree_26)|n121_tree_26;
    assign n122_tree_26 = a_in[20]|b_in[20];

    assign n121_tree_26 = a_in[20]&b_in[20];
    assign n123_tree_26 = (n126_tree_26&n125_tree_26)|n124_tree_26;
    assign n125_tree_26 = a_in[19]|b_in[19];

    assign n124_tree_26 = a_in[19]&b_in[19];
    assign n126_tree_26 = (n129_tree_26&n128_tree_26)|n127_tree_26;
    assign n128_tree_26 = a_in[18]|b_in[18];

    assign n127_tree_26 = a_in[18]&b_in[18];
    assign n129_tree_26 = (n132_tree_26&n131_tree_26)|n130_tree_26;
    assign n131_tree_26 = a_in[17]|b_in[17];

    assign n130_tree_26 = a_in[17]&b_in[17];
    assign n132_tree_26 = (n135_tree_26&n134_tree_26)|n133_tree_26;
    assign n134_tree_26 = a_in[16]|b_in[16];

    assign n133_tree_26 = a_in[16]&b_in[16];
    assign n135_tree_26 = (n138_tree_26&n137_tree_26)|n136_tree_26;
    assign n137_tree_26 = a_in[15]|b_in[15];

    assign n136_tree_26 = a_in[15]&b_in[15];
    assign n138_tree_26 = (n141_tree_26&n140_tree_26)|n139_tree_26;
    assign n140_tree_26 = a_in[14]|b_in[14];

    assign n139_tree_26 = a_in[14]&b_in[14];
    assign n141_tree_26 = (n144_tree_26&n143_tree_26)|n142_tree_26;
    assign n143_tree_26 = a_in[13]|b_in[13];

    assign n142_tree_26 = a_in[13]&b_in[13];
    assign n144_tree_26 = (n147_tree_26&n146_tree_26)|n145_tree_26;
    assign n146_tree_26 = a_in[12]|b_in[12];

    assign n145_tree_26 = a_in[12]&b_in[12];
    assign n147_tree_26 = (n150_tree_26&n149_tree_26)|n148_tree_26;
    assign n149_tree_26 = a_in[11]|b_in[11];

    assign n148_tree_26 = a_in[11]&b_in[11];
    assign n150_tree_26 = (n153_tree_26&n152_tree_26)|n151_tree_26;
    assign n152_tree_26 = a_in[10]|b_in[10];

    assign n151_tree_26 = a_in[10]&b_in[10];
    assign n153_tree_26 = (n156_tree_26&n155_tree_26)|n154_tree_26;
    assign n155_tree_26 = a_in[9]|b_in[9];

    assign n154_tree_26 = a_in[9]&b_in[9];
    assign n156_tree_26 = (n159_tree_26&n158_tree_26)|n157_tree_26;
    assign n158_tree_26 = a_in[8]|b_in[8];

    assign n157_tree_26 = a_in[8]&b_in[8];
    assign n159_tree_26 = (n162_tree_26&n161_tree_26)|n160_tree_26;
    assign n161_tree_26 = a_in[7]|b_in[7];

    assign n160_tree_26 = a_in[7]&b_in[7];
    assign n162_tree_26 = (n165_tree_26&n164_tree_26)|n163_tree_26;
    assign n164_tree_26 = a_in[6]|b_in[6];

    assign n163_tree_26 = a_in[6]&b_in[6];
    assign n165_tree_26 = (n168_tree_26&n167_tree_26)|n166_tree_26;
    assign n167_tree_26 = a_in[5]|b_in[5];

    assign n166_tree_26 = a_in[5]&b_in[5];
    assign n168_tree_26 = (n171_tree_26&n170_tree_26)|n169_tree_26;
    assign n170_tree_26 = a_in[4]|b_in[4];

    assign n169_tree_26 = a_in[4]&b_in[4];
    assign n171_tree_26 = (n174_tree_26&n173_tree_26)|n172_tree_26;
    assign n173_tree_26 = a_in[3]|b_in[3];

    assign n172_tree_26 = a_in[3]&b_in[3];
    assign n174_tree_26 = (n177_tree_26&n176_tree_26)|n175_tree_26;
    assign n176_tree_26 = a_in[2]|b_in[2];

    assign n175_tree_26 = a_in[2]&b_in[2];
    assign n177_tree_26 = (n180_tree_26&n179_tree_26)|n178_tree_26;
    assign n179_tree_26 = a_in[1]|b_in[1];

    assign n178_tree_26 = a_in[1]&b_in[1];
    assign n180_tree_26 = a_in[0]&b_in[0];

// adder_forest tree_25
	wire n100_tree_25, n101_tree_25, n102_tree_25, n103_tree_25, n104_tree_25, n105_tree_25, n106_tree_25, n107_tree_25, n108_tree_25, n109_tree_25, n110_tree_25, n111_tree_25, n112_tree_25, n113_tree_25, n114_tree_25, n115_tree_25, n116_tree_25, n117_tree_25, n118_tree_25, n119_tree_25, n120_tree_25, n121_tree_25, n122_tree_25, n123_tree_25, n124_tree_25, n125_tree_25, n126_tree_25, n127_tree_25, n128_tree_25, n129_tree_25, n130_tree_25, n131_tree_25, n132_tree_25, n133_tree_25, n134_tree_25, n135_tree_25, n136_tree_25, n137_tree_25, n138_tree_25, n139_tree_25, n140_tree_25, n141_tree_25, n142_tree_25, n143_tree_25, n144_tree_25, n145_tree_25, n146_tree_25, n147_tree_25, n148_tree_25, n149_tree_25, n150_tree_25, n151_tree_25, n152_tree_25, n153_tree_25, n154_tree_25, n155_tree_25, n156_tree_25, n157_tree_25, n158_tree_25, n159_tree_25, n160_tree_25, n161_tree_25, n162_tree_25, n163_tree_25, n164_tree_25, n165_tree_25, n166_tree_25, n167_tree_25, n168_tree_25, n169_tree_25, n170_tree_25, n171_tree_25, n172_tree_25, n173_tree_25;
    assign sum[25] = n101_tree_25^n100_tree_25;
    assign n100_tree_25 = a_in[25]^b_in[25];
    assign n101_tree_25 = (n104_tree_25&n103_tree_25)|n102_tree_25;
    assign n103_tree_25 = a_in[24]|b_in[24];

    assign n102_tree_25 = a_in[24]&b_in[24];
    assign n104_tree_25 = (n107_tree_25&n106_tree_25)|n105_tree_25;
    assign n106_tree_25 = a_in[23]|b_in[23];

    assign n105_tree_25 = a_in[23]&b_in[23];
    assign n107_tree_25 = (n110_tree_25&n109_tree_25)|n108_tree_25;
    assign n109_tree_25 = a_in[22]|b_in[22];

    assign n108_tree_25 = a_in[22]&b_in[22];
    assign n110_tree_25 = (n113_tree_25&n112_tree_25)|n111_tree_25;
    assign n112_tree_25 = a_in[21]|b_in[21];

    assign n111_tree_25 = a_in[21]&b_in[21];
    assign n113_tree_25 = (n116_tree_25&n115_tree_25)|n114_tree_25;
    assign n115_tree_25 = a_in[20]|b_in[20];

    assign n114_tree_25 = a_in[20]&b_in[20];
    assign n116_tree_25 = (n119_tree_25&n118_tree_25)|n117_tree_25;
    assign n118_tree_25 = a_in[19]|b_in[19];

    assign n117_tree_25 = a_in[19]&b_in[19];
    assign n119_tree_25 = (n122_tree_25&n121_tree_25)|n120_tree_25;
    assign n121_tree_25 = a_in[18]|b_in[18];

    assign n120_tree_25 = a_in[18]&b_in[18];
    assign n122_tree_25 = (n125_tree_25&n124_tree_25)|n123_tree_25;
    assign n124_tree_25 = a_in[17]|b_in[17];

    assign n123_tree_25 = a_in[17]&b_in[17];
    assign n125_tree_25 = (n128_tree_25&n127_tree_25)|n126_tree_25;
    assign n127_tree_25 = a_in[16]|b_in[16];

    assign n126_tree_25 = a_in[16]&b_in[16];
    assign n128_tree_25 = (n131_tree_25&n130_tree_25)|n129_tree_25;
    assign n130_tree_25 = a_in[15]|b_in[15];

    assign n129_tree_25 = a_in[15]&b_in[15];
    assign n131_tree_25 = (n134_tree_25&n133_tree_25)|n132_tree_25;
    assign n133_tree_25 = a_in[14]|b_in[14];

    assign n132_tree_25 = a_in[14]&b_in[14];
    assign n134_tree_25 = (n137_tree_25&n136_tree_25)|n135_tree_25;
    assign n136_tree_25 = a_in[13]|b_in[13];

    assign n135_tree_25 = a_in[13]&b_in[13];
    assign n137_tree_25 = (n140_tree_25&n139_tree_25)|n138_tree_25;
    assign n139_tree_25 = a_in[12]|b_in[12];

    assign n138_tree_25 = a_in[12]&b_in[12];
    assign n140_tree_25 = (n143_tree_25&n142_tree_25)|n141_tree_25;
    assign n142_tree_25 = a_in[11]|b_in[11];

    assign n141_tree_25 = a_in[11]&b_in[11];
    assign n143_tree_25 = (n146_tree_25&n145_tree_25)|n144_tree_25;
    assign n145_tree_25 = a_in[10]|b_in[10];

    assign n144_tree_25 = a_in[10]&b_in[10];
    assign n146_tree_25 = (n149_tree_25&n148_tree_25)|n147_tree_25;
    assign n148_tree_25 = a_in[9]|b_in[9];

    assign n147_tree_25 = a_in[9]&b_in[9];
    assign n149_tree_25 = (n152_tree_25&n151_tree_25)|n150_tree_25;
    assign n151_tree_25 = a_in[8]|b_in[8];

    assign n150_tree_25 = a_in[8]&b_in[8];
    assign n152_tree_25 = (n155_tree_25&n154_tree_25)|n153_tree_25;
    assign n154_tree_25 = a_in[7]|b_in[7];

    assign n153_tree_25 = a_in[7]&b_in[7];
    assign n155_tree_25 = (n158_tree_25&n157_tree_25)|n156_tree_25;
    assign n157_tree_25 = a_in[6]|b_in[6];

    assign n156_tree_25 = a_in[6]&b_in[6];
    assign n158_tree_25 = (n161_tree_25&n160_tree_25)|n159_tree_25;
    assign n160_tree_25 = a_in[5]|b_in[5];

    assign n159_tree_25 = a_in[5]&b_in[5];
    assign n161_tree_25 = (n164_tree_25&n163_tree_25)|n162_tree_25;
    assign n163_tree_25 = a_in[4]|b_in[4];

    assign n162_tree_25 = a_in[4]&b_in[4];
    assign n164_tree_25 = (n167_tree_25&n166_tree_25)|n165_tree_25;
    assign n166_tree_25 = a_in[3]|b_in[3];

    assign n165_tree_25 = a_in[3]&b_in[3];
    assign n167_tree_25 = (n170_tree_25&n169_tree_25)|n168_tree_25;
    assign n169_tree_25 = a_in[2]|b_in[2];

    assign n168_tree_25 = a_in[2]&b_in[2];
    assign n170_tree_25 = (n173_tree_25&n172_tree_25)|n171_tree_25;
    assign n172_tree_25 = a_in[1]|b_in[1];

    assign n171_tree_25 = a_in[1]&b_in[1];
    assign n173_tree_25 = a_in[0]&b_in[0];

// adder_forest tree_24
	wire n96_tree_24, n97_tree_24, n98_tree_24, n99_tree_24, n100_tree_24, n101_tree_24, n102_tree_24, n103_tree_24, n104_tree_24, n105_tree_24, n106_tree_24, n107_tree_24, n108_tree_24, n109_tree_24, n110_tree_24, n111_tree_24, n112_tree_24, n113_tree_24, n114_tree_24, n115_tree_24, n116_tree_24, n117_tree_24, n118_tree_24, n119_tree_24, n120_tree_24, n121_tree_24, n122_tree_24, n123_tree_24, n124_tree_24, n125_tree_24, n126_tree_24, n127_tree_24, n128_tree_24, n129_tree_24, n130_tree_24, n131_tree_24, n132_tree_24, n133_tree_24, n134_tree_24, n135_tree_24, n136_tree_24, n137_tree_24, n138_tree_24, n139_tree_24, n140_tree_24, n141_tree_24, n142_tree_24, n143_tree_24, n144_tree_24, n145_tree_24, n146_tree_24, n147_tree_24, n148_tree_24, n149_tree_24, n150_tree_24, n151_tree_24, n152_tree_24, n153_tree_24, n154_tree_24, n155_tree_24, n156_tree_24, n157_tree_24, n158_tree_24, n159_tree_24, n160_tree_24, n161_tree_24, n162_tree_24, n163_tree_24, n164_tree_24, n165_tree_24, n166_tree_24;
    assign sum[24] = n97_tree_24^n96_tree_24;
    assign n96_tree_24 = a_in[24]^b_in[24];
    assign n97_tree_24 = (n100_tree_24&n99_tree_24)|n98_tree_24;
    assign n99_tree_24 = a_in[23]|b_in[23];

    assign n98_tree_24 = a_in[23]&b_in[23];
    assign n100_tree_24 = (n103_tree_24&n102_tree_24)|n101_tree_24;
    assign n102_tree_24 = a_in[22]|b_in[22];

    assign n101_tree_24 = a_in[22]&b_in[22];
    assign n103_tree_24 = (n106_tree_24&n105_tree_24)|n104_tree_24;
    assign n105_tree_24 = a_in[21]|b_in[21];

    assign n104_tree_24 = a_in[21]&b_in[21];
    assign n106_tree_24 = (n109_tree_24&n108_tree_24)|n107_tree_24;
    assign n108_tree_24 = a_in[20]|b_in[20];

    assign n107_tree_24 = a_in[20]&b_in[20];
    assign n109_tree_24 = (n112_tree_24&n111_tree_24)|n110_tree_24;
    assign n111_tree_24 = a_in[19]|b_in[19];

    assign n110_tree_24 = a_in[19]&b_in[19];
    assign n112_tree_24 = (n115_tree_24&n114_tree_24)|n113_tree_24;
    assign n114_tree_24 = a_in[18]|b_in[18];

    assign n113_tree_24 = a_in[18]&b_in[18];
    assign n115_tree_24 = (n118_tree_24&n117_tree_24)|n116_tree_24;
    assign n117_tree_24 = a_in[17]|b_in[17];

    assign n116_tree_24 = a_in[17]&b_in[17];
    assign n118_tree_24 = (n121_tree_24&n120_tree_24)|n119_tree_24;
    assign n120_tree_24 = a_in[16]|b_in[16];

    assign n119_tree_24 = a_in[16]&b_in[16];
    assign n121_tree_24 = (n124_tree_24&n123_tree_24)|n122_tree_24;
    assign n123_tree_24 = a_in[15]|b_in[15];

    assign n122_tree_24 = a_in[15]&b_in[15];
    assign n124_tree_24 = (n127_tree_24&n126_tree_24)|n125_tree_24;
    assign n126_tree_24 = a_in[14]|b_in[14];

    assign n125_tree_24 = a_in[14]&b_in[14];
    assign n127_tree_24 = (n130_tree_24&n129_tree_24)|n128_tree_24;
    assign n129_tree_24 = a_in[13]|b_in[13];

    assign n128_tree_24 = a_in[13]&b_in[13];
    assign n130_tree_24 = (n133_tree_24&n132_tree_24)|n131_tree_24;
    assign n132_tree_24 = a_in[12]|b_in[12];

    assign n131_tree_24 = a_in[12]&b_in[12];
    assign n133_tree_24 = (n136_tree_24&n135_tree_24)|n134_tree_24;
    assign n135_tree_24 = a_in[11]|b_in[11];

    assign n134_tree_24 = a_in[11]&b_in[11];
    assign n136_tree_24 = (n139_tree_24&n138_tree_24)|n137_tree_24;
    assign n138_tree_24 = a_in[10]|b_in[10];

    assign n137_tree_24 = a_in[10]&b_in[10];
    assign n139_tree_24 = (n142_tree_24&n141_tree_24)|n140_tree_24;
    assign n141_tree_24 = a_in[9]|b_in[9];

    assign n140_tree_24 = a_in[9]&b_in[9];
    assign n142_tree_24 = (n145_tree_24&n144_tree_24)|n143_tree_24;
    assign n144_tree_24 = a_in[8]|b_in[8];

    assign n143_tree_24 = a_in[8]&b_in[8];
    assign n145_tree_24 = (n148_tree_24&n147_tree_24)|n146_tree_24;
    assign n147_tree_24 = a_in[7]|b_in[7];

    assign n146_tree_24 = a_in[7]&b_in[7];
    assign n148_tree_24 = (n151_tree_24&n150_tree_24)|n149_tree_24;
    assign n150_tree_24 = a_in[6]|b_in[6];

    assign n149_tree_24 = a_in[6]&b_in[6];
    assign n151_tree_24 = (n154_tree_24&n153_tree_24)|n152_tree_24;
    assign n153_tree_24 = a_in[5]|b_in[5];

    assign n152_tree_24 = a_in[5]&b_in[5];
    assign n154_tree_24 = (n157_tree_24&n156_tree_24)|n155_tree_24;
    assign n156_tree_24 = a_in[4]|b_in[4];

    assign n155_tree_24 = a_in[4]&b_in[4];
    assign n157_tree_24 = (n160_tree_24&n159_tree_24)|n158_tree_24;
    assign n159_tree_24 = a_in[3]|b_in[3];

    assign n158_tree_24 = a_in[3]&b_in[3];
    assign n160_tree_24 = (n163_tree_24&n162_tree_24)|n161_tree_24;
    assign n162_tree_24 = a_in[2]|b_in[2];

    assign n161_tree_24 = a_in[2]&b_in[2];
    assign n163_tree_24 = (n166_tree_24&n165_tree_24)|n164_tree_24;
    assign n165_tree_24 = a_in[1]|b_in[1];

    assign n164_tree_24 = a_in[1]&b_in[1];
    assign n166_tree_24 = a_in[0]&b_in[0];

// adder_forest tree_23
	wire n92_tree_23, n93_tree_23, n94_tree_23, n95_tree_23, n96_tree_23, n97_tree_23, n98_tree_23, n99_tree_23, n100_tree_23, n101_tree_23, n102_tree_23, n103_tree_23, n104_tree_23, n105_tree_23, n106_tree_23, n107_tree_23, n108_tree_23, n109_tree_23, n110_tree_23, n111_tree_23, n112_tree_23, n113_tree_23, n114_tree_23, n115_tree_23, n116_tree_23, n117_tree_23, n118_tree_23, n119_tree_23, n120_tree_23, n121_tree_23, n122_tree_23, n123_tree_23, n124_tree_23, n125_tree_23, n126_tree_23, n127_tree_23, n128_tree_23, n129_tree_23, n130_tree_23, n131_tree_23, n132_tree_23, n133_tree_23, n134_tree_23, n135_tree_23, n136_tree_23, n137_tree_23, n138_tree_23, n139_tree_23, n140_tree_23, n141_tree_23, n142_tree_23, n143_tree_23, n144_tree_23, n145_tree_23, n146_tree_23, n147_tree_23, n148_tree_23, n149_tree_23, n150_tree_23, n151_tree_23, n152_tree_23, n153_tree_23, n154_tree_23, n155_tree_23, n156_tree_23, n157_tree_23, n158_tree_23, n159_tree_23;
    assign sum[23] = n93_tree_23^n92_tree_23;
    assign n92_tree_23 = a_in[23]^b_in[23];
    assign n93_tree_23 = (n96_tree_23&n95_tree_23)|n94_tree_23;
    assign n95_tree_23 = a_in[22]|b_in[22];

    assign n94_tree_23 = a_in[22]&b_in[22];
    assign n96_tree_23 = (n99_tree_23&n98_tree_23)|n97_tree_23;
    assign n98_tree_23 = a_in[21]|b_in[21];

    assign n97_tree_23 = a_in[21]&b_in[21];
    assign n99_tree_23 = (n102_tree_23&n101_tree_23)|n100_tree_23;
    assign n101_tree_23 = a_in[20]|b_in[20];

    assign n100_tree_23 = a_in[20]&b_in[20];
    assign n102_tree_23 = (n105_tree_23&n104_tree_23)|n103_tree_23;
    assign n104_tree_23 = a_in[19]|b_in[19];

    assign n103_tree_23 = a_in[19]&b_in[19];
    assign n105_tree_23 = (n108_tree_23&n107_tree_23)|n106_tree_23;
    assign n107_tree_23 = a_in[18]|b_in[18];

    assign n106_tree_23 = a_in[18]&b_in[18];
    assign n108_tree_23 = (n111_tree_23&n110_tree_23)|n109_tree_23;
    assign n110_tree_23 = a_in[17]|b_in[17];

    assign n109_tree_23 = a_in[17]&b_in[17];
    assign n111_tree_23 = (n114_tree_23&n113_tree_23)|n112_tree_23;
    assign n113_tree_23 = a_in[16]|b_in[16];

    assign n112_tree_23 = a_in[16]&b_in[16];
    assign n114_tree_23 = (n117_tree_23&n116_tree_23)|n115_tree_23;
    assign n116_tree_23 = a_in[15]|b_in[15];

    assign n115_tree_23 = a_in[15]&b_in[15];
    assign n117_tree_23 = (n120_tree_23&n119_tree_23)|n118_tree_23;
    assign n119_tree_23 = a_in[14]|b_in[14];

    assign n118_tree_23 = a_in[14]&b_in[14];
    assign n120_tree_23 = (n123_tree_23&n122_tree_23)|n121_tree_23;
    assign n122_tree_23 = a_in[13]|b_in[13];

    assign n121_tree_23 = a_in[13]&b_in[13];
    assign n123_tree_23 = (n126_tree_23&n125_tree_23)|n124_tree_23;
    assign n125_tree_23 = a_in[12]|b_in[12];

    assign n124_tree_23 = a_in[12]&b_in[12];
    assign n126_tree_23 = (n129_tree_23&n128_tree_23)|n127_tree_23;
    assign n128_tree_23 = a_in[11]|b_in[11];

    assign n127_tree_23 = a_in[11]&b_in[11];
    assign n129_tree_23 = (n132_tree_23&n131_tree_23)|n130_tree_23;
    assign n131_tree_23 = a_in[10]|b_in[10];

    assign n130_tree_23 = a_in[10]&b_in[10];
    assign n132_tree_23 = (n135_tree_23&n134_tree_23)|n133_tree_23;
    assign n134_tree_23 = a_in[9]|b_in[9];

    assign n133_tree_23 = a_in[9]&b_in[9];
    assign n135_tree_23 = (n138_tree_23&n137_tree_23)|n136_tree_23;
    assign n137_tree_23 = a_in[8]|b_in[8];

    assign n136_tree_23 = a_in[8]&b_in[8];
    assign n138_tree_23 = (n141_tree_23&n140_tree_23)|n139_tree_23;
    assign n140_tree_23 = a_in[7]|b_in[7];

    assign n139_tree_23 = a_in[7]&b_in[7];
    assign n141_tree_23 = (n144_tree_23&n143_tree_23)|n142_tree_23;
    assign n143_tree_23 = a_in[6]|b_in[6];

    assign n142_tree_23 = a_in[6]&b_in[6];
    assign n144_tree_23 = (n147_tree_23&n146_tree_23)|n145_tree_23;
    assign n146_tree_23 = a_in[5]|b_in[5];

    assign n145_tree_23 = a_in[5]&b_in[5];
    assign n147_tree_23 = (n150_tree_23&n149_tree_23)|n148_tree_23;
    assign n149_tree_23 = a_in[4]|b_in[4];

    assign n148_tree_23 = a_in[4]&b_in[4];
    assign n150_tree_23 = (n153_tree_23&n152_tree_23)|n151_tree_23;
    assign n152_tree_23 = a_in[3]|b_in[3];

    assign n151_tree_23 = a_in[3]&b_in[3];
    assign n153_tree_23 = (n156_tree_23&n155_tree_23)|n154_tree_23;
    assign n155_tree_23 = a_in[2]|b_in[2];

    assign n154_tree_23 = a_in[2]&b_in[2];
    assign n156_tree_23 = (n159_tree_23&n158_tree_23)|n157_tree_23;
    assign n158_tree_23 = a_in[1]|b_in[1];

    assign n157_tree_23 = a_in[1]&b_in[1];
    assign n159_tree_23 = a_in[0]&b_in[0];

// adder_forest tree_22
	wire n88_tree_22, n89_tree_22, n90_tree_22, n91_tree_22, n92_tree_22, n93_tree_22, n94_tree_22, n95_tree_22, n96_tree_22, n97_tree_22, n98_tree_22, n99_tree_22, n100_tree_22, n101_tree_22, n102_tree_22, n103_tree_22, n104_tree_22, n105_tree_22, n106_tree_22, n107_tree_22, n108_tree_22, n109_tree_22, n110_tree_22, n111_tree_22, n112_tree_22, n113_tree_22, n114_tree_22, n115_tree_22, n116_tree_22, n117_tree_22, n118_tree_22, n119_tree_22, n120_tree_22, n121_tree_22, n122_tree_22, n123_tree_22, n124_tree_22, n125_tree_22, n126_tree_22, n127_tree_22, n128_tree_22, n129_tree_22, n130_tree_22, n131_tree_22, n132_tree_22, n133_tree_22, n134_tree_22, n135_tree_22, n136_tree_22, n137_tree_22, n138_tree_22, n139_tree_22, n140_tree_22, n141_tree_22, n142_tree_22, n143_tree_22, n144_tree_22, n145_tree_22, n146_tree_22, n147_tree_22, n148_tree_22, n149_tree_22, n150_tree_22, n151_tree_22, n152_tree_22;
    assign sum[22] = n89_tree_22^n88_tree_22;
    assign n88_tree_22 = a_in[22]^b_in[22];
    assign n89_tree_22 = (n92_tree_22&n91_tree_22)|n90_tree_22;
    assign n91_tree_22 = a_in[21]|b_in[21];

    assign n90_tree_22 = a_in[21]&b_in[21];
    assign n92_tree_22 = (n95_tree_22&n94_tree_22)|n93_tree_22;
    assign n94_tree_22 = a_in[20]|b_in[20];

    assign n93_tree_22 = a_in[20]&b_in[20];
    assign n95_tree_22 = (n98_tree_22&n97_tree_22)|n96_tree_22;
    assign n97_tree_22 = a_in[19]|b_in[19];

    assign n96_tree_22 = a_in[19]&b_in[19];
    assign n98_tree_22 = (n101_tree_22&n100_tree_22)|n99_tree_22;
    assign n100_tree_22 = a_in[18]|b_in[18];

    assign n99_tree_22 = a_in[18]&b_in[18];
    assign n101_tree_22 = (n104_tree_22&n103_tree_22)|n102_tree_22;
    assign n103_tree_22 = a_in[17]|b_in[17];

    assign n102_tree_22 = a_in[17]&b_in[17];
    assign n104_tree_22 = (n107_tree_22&n106_tree_22)|n105_tree_22;
    assign n106_tree_22 = a_in[16]|b_in[16];

    assign n105_tree_22 = a_in[16]&b_in[16];
    assign n107_tree_22 = (n110_tree_22&n109_tree_22)|n108_tree_22;
    assign n109_tree_22 = a_in[15]|b_in[15];

    assign n108_tree_22 = a_in[15]&b_in[15];
    assign n110_tree_22 = (n113_tree_22&n112_tree_22)|n111_tree_22;
    assign n112_tree_22 = a_in[14]|b_in[14];

    assign n111_tree_22 = a_in[14]&b_in[14];
    assign n113_tree_22 = (n116_tree_22&n115_tree_22)|n114_tree_22;
    assign n115_tree_22 = a_in[13]|b_in[13];

    assign n114_tree_22 = a_in[13]&b_in[13];
    assign n116_tree_22 = (n119_tree_22&n118_tree_22)|n117_tree_22;
    assign n118_tree_22 = a_in[12]|b_in[12];

    assign n117_tree_22 = a_in[12]&b_in[12];
    assign n119_tree_22 = (n122_tree_22&n121_tree_22)|n120_tree_22;
    assign n121_tree_22 = a_in[11]|b_in[11];

    assign n120_tree_22 = a_in[11]&b_in[11];
    assign n122_tree_22 = (n125_tree_22&n124_tree_22)|n123_tree_22;
    assign n124_tree_22 = a_in[10]|b_in[10];

    assign n123_tree_22 = a_in[10]&b_in[10];
    assign n125_tree_22 = (n128_tree_22&n127_tree_22)|n126_tree_22;
    assign n127_tree_22 = a_in[9]|b_in[9];

    assign n126_tree_22 = a_in[9]&b_in[9];
    assign n128_tree_22 = (n131_tree_22&n130_tree_22)|n129_tree_22;
    assign n130_tree_22 = a_in[8]|b_in[8];

    assign n129_tree_22 = a_in[8]&b_in[8];
    assign n131_tree_22 = (n134_tree_22&n133_tree_22)|n132_tree_22;
    assign n133_tree_22 = a_in[7]|b_in[7];

    assign n132_tree_22 = a_in[7]&b_in[7];
    assign n134_tree_22 = (n137_tree_22&n136_tree_22)|n135_tree_22;
    assign n136_tree_22 = a_in[6]|b_in[6];

    assign n135_tree_22 = a_in[6]&b_in[6];
    assign n137_tree_22 = (n140_tree_22&n139_tree_22)|n138_tree_22;
    assign n139_tree_22 = a_in[5]|b_in[5];

    assign n138_tree_22 = a_in[5]&b_in[5];
    assign n140_tree_22 = (n143_tree_22&n142_tree_22)|n141_tree_22;
    assign n142_tree_22 = a_in[4]|b_in[4];

    assign n141_tree_22 = a_in[4]&b_in[4];
    assign n143_tree_22 = (n146_tree_22&n145_tree_22)|n144_tree_22;
    assign n145_tree_22 = a_in[3]|b_in[3];

    assign n144_tree_22 = a_in[3]&b_in[3];
    assign n146_tree_22 = (n149_tree_22&n148_tree_22)|n147_tree_22;
    assign n148_tree_22 = a_in[2]|b_in[2];

    assign n147_tree_22 = a_in[2]&b_in[2];
    assign n149_tree_22 = (n152_tree_22&n151_tree_22)|n150_tree_22;
    assign n151_tree_22 = a_in[1]|b_in[1];

    assign n150_tree_22 = a_in[1]&b_in[1];
    assign n152_tree_22 = a_in[0]&b_in[0];

// adder_forest tree_21
	wire n84_tree_21, n85_tree_21, n86_tree_21, n87_tree_21, n88_tree_21, n89_tree_21, n90_tree_21, n91_tree_21, n92_tree_21, n93_tree_21, n94_tree_21, n95_tree_21, n96_tree_21, n97_tree_21, n98_tree_21, n99_tree_21, n100_tree_21, n101_tree_21, n102_tree_21, n103_tree_21, n104_tree_21, n105_tree_21, n106_tree_21, n107_tree_21, n108_tree_21, n109_tree_21, n110_tree_21, n111_tree_21, n112_tree_21, n113_tree_21, n114_tree_21, n115_tree_21, n116_tree_21, n117_tree_21, n118_tree_21, n119_tree_21, n120_tree_21, n121_tree_21, n122_tree_21, n123_tree_21, n124_tree_21, n125_tree_21, n126_tree_21, n127_tree_21, n128_tree_21, n129_tree_21, n130_tree_21, n131_tree_21, n132_tree_21, n133_tree_21, n134_tree_21, n135_tree_21, n136_tree_21, n137_tree_21, n138_tree_21, n139_tree_21, n140_tree_21, n141_tree_21, n142_tree_21, n143_tree_21, n144_tree_21, n145_tree_21;
    assign sum[21] = n85_tree_21^n84_tree_21;
    assign n84_tree_21 = a_in[21]^b_in[21];
    assign n85_tree_21 = (n88_tree_21&n87_tree_21)|n86_tree_21;
    assign n87_tree_21 = a_in[20]|b_in[20];

    assign n86_tree_21 = a_in[20]&b_in[20];
    assign n88_tree_21 = (n91_tree_21&n90_tree_21)|n89_tree_21;
    assign n90_tree_21 = a_in[19]|b_in[19];

    assign n89_tree_21 = a_in[19]&b_in[19];
    assign n91_tree_21 = (n94_tree_21&n93_tree_21)|n92_tree_21;
    assign n93_tree_21 = a_in[18]|b_in[18];

    assign n92_tree_21 = a_in[18]&b_in[18];
    assign n94_tree_21 = (n97_tree_21&n96_tree_21)|n95_tree_21;
    assign n96_tree_21 = a_in[17]|b_in[17];

    assign n95_tree_21 = a_in[17]&b_in[17];
    assign n97_tree_21 = (n100_tree_21&n99_tree_21)|n98_tree_21;
    assign n99_tree_21 = a_in[16]|b_in[16];

    assign n98_tree_21 = a_in[16]&b_in[16];
    assign n100_tree_21 = (n103_tree_21&n102_tree_21)|n101_tree_21;
    assign n102_tree_21 = a_in[15]|b_in[15];

    assign n101_tree_21 = a_in[15]&b_in[15];
    assign n103_tree_21 = (n106_tree_21&n105_tree_21)|n104_tree_21;
    assign n105_tree_21 = a_in[14]|b_in[14];

    assign n104_tree_21 = a_in[14]&b_in[14];
    assign n106_tree_21 = (n109_tree_21&n108_tree_21)|n107_tree_21;
    assign n108_tree_21 = a_in[13]|b_in[13];

    assign n107_tree_21 = a_in[13]&b_in[13];
    assign n109_tree_21 = (n112_tree_21&n111_tree_21)|n110_tree_21;
    assign n111_tree_21 = a_in[12]|b_in[12];

    assign n110_tree_21 = a_in[12]&b_in[12];
    assign n112_tree_21 = (n115_tree_21&n114_tree_21)|n113_tree_21;
    assign n114_tree_21 = a_in[11]|b_in[11];

    assign n113_tree_21 = a_in[11]&b_in[11];
    assign n115_tree_21 = (n118_tree_21&n117_tree_21)|n116_tree_21;
    assign n117_tree_21 = a_in[10]|b_in[10];

    assign n116_tree_21 = a_in[10]&b_in[10];
    assign n118_tree_21 = (n121_tree_21&n120_tree_21)|n119_tree_21;
    assign n120_tree_21 = a_in[9]|b_in[9];

    assign n119_tree_21 = a_in[9]&b_in[9];
    assign n121_tree_21 = (n124_tree_21&n123_tree_21)|n122_tree_21;
    assign n123_tree_21 = a_in[8]|b_in[8];

    assign n122_tree_21 = a_in[8]&b_in[8];
    assign n124_tree_21 = (n127_tree_21&n126_tree_21)|n125_tree_21;
    assign n126_tree_21 = a_in[7]|b_in[7];

    assign n125_tree_21 = a_in[7]&b_in[7];
    assign n127_tree_21 = (n130_tree_21&n129_tree_21)|n128_tree_21;
    assign n129_tree_21 = a_in[6]|b_in[6];

    assign n128_tree_21 = a_in[6]&b_in[6];
    assign n130_tree_21 = (n133_tree_21&n132_tree_21)|n131_tree_21;
    assign n132_tree_21 = a_in[5]|b_in[5];

    assign n131_tree_21 = a_in[5]&b_in[5];
    assign n133_tree_21 = (n136_tree_21&n135_tree_21)|n134_tree_21;
    assign n135_tree_21 = a_in[4]|b_in[4];

    assign n134_tree_21 = a_in[4]&b_in[4];
    assign n136_tree_21 = (n139_tree_21&n138_tree_21)|n137_tree_21;
    assign n138_tree_21 = a_in[3]|b_in[3];

    assign n137_tree_21 = a_in[3]&b_in[3];
    assign n139_tree_21 = (n142_tree_21&n141_tree_21)|n140_tree_21;
    assign n141_tree_21 = a_in[2]|b_in[2];

    assign n140_tree_21 = a_in[2]&b_in[2];
    assign n142_tree_21 = (n145_tree_21&n144_tree_21)|n143_tree_21;
    assign n144_tree_21 = a_in[1]|b_in[1];

    assign n143_tree_21 = a_in[1]&b_in[1];
    assign n145_tree_21 = a_in[0]&b_in[0];

// adder_forest tree_20
	wire n80_tree_20, n81_tree_20, n82_tree_20, n83_tree_20, n84_tree_20, n85_tree_20, n86_tree_20, n87_tree_20, n88_tree_20, n89_tree_20, n90_tree_20, n91_tree_20, n92_tree_20, n93_tree_20, n94_tree_20, n95_tree_20, n96_tree_20, n97_tree_20, n98_tree_20, n99_tree_20, n100_tree_20, n101_tree_20, n102_tree_20, n103_tree_20, n104_tree_20, n105_tree_20, n106_tree_20, n107_tree_20, n108_tree_20, n109_tree_20, n110_tree_20, n111_tree_20, n112_tree_20, n113_tree_20, n114_tree_20, n115_tree_20, n116_tree_20, n117_tree_20, n118_tree_20, n119_tree_20, n120_tree_20, n121_tree_20, n122_tree_20, n123_tree_20, n124_tree_20, n125_tree_20, n126_tree_20, n127_tree_20, n128_tree_20, n129_tree_20, n130_tree_20, n131_tree_20, n132_tree_20, n133_tree_20, n134_tree_20, n135_tree_20, n136_tree_20, n137_tree_20, n138_tree_20;
    assign sum[20] = n81_tree_20^n80_tree_20;
    assign n80_tree_20 = a_in[20]^b_in[20];
    assign n81_tree_20 = (n84_tree_20&n83_tree_20)|n82_tree_20;
    assign n83_tree_20 = a_in[19]|b_in[19];

    assign n82_tree_20 = a_in[19]&b_in[19];
    assign n84_tree_20 = (n87_tree_20&n86_tree_20)|n85_tree_20;
    assign n86_tree_20 = a_in[18]|b_in[18];

    assign n85_tree_20 = a_in[18]&b_in[18];
    assign n87_tree_20 = (n90_tree_20&n89_tree_20)|n88_tree_20;
    assign n89_tree_20 = a_in[17]|b_in[17];

    assign n88_tree_20 = a_in[17]&b_in[17];
    assign n90_tree_20 = (n93_tree_20&n92_tree_20)|n91_tree_20;
    assign n92_tree_20 = a_in[16]|b_in[16];

    assign n91_tree_20 = a_in[16]&b_in[16];
    assign n93_tree_20 = (n96_tree_20&n95_tree_20)|n94_tree_20;
    assign n95_tree_20 = a_in[15]|b_in[15];

    assign n94_tree_20 = a_in[15]&b_in[15];
    assign n96_tree_20 = (n99_tree_20&n98_tree_20)|n97_tree_20;
    assign n98_tree_20 = a_in[14]|b_in[14];

    assign n97_tree_20 = a_in[14]&b_in[14];
    assign n99_tree_20 = (n102_tree_20&n101_tree_20)|n100_tree_20;
    assign n101_tree_20 = a_in[13]|b_in[13];

    assign n100_tree_20 = a_in[13]&b_in[13];
    assign n102_tree_20 = (n105_tree_20&n104_tree_20)|n103_tree_20;
    assign n104_tree_20 = a_in[12]|b_in[12];

    assign n103_tree_20 = a_in[12]&b_in[12];
    assign n105_tree_20 = (n108_tree_20&n107_tree_20)|n106_tree_20;
    assign n107_tree_20 = a_in[11]|b_in[11];

    assign n106_tree_20 = a_in[11]&b_in[11];
    assign n108_tree_20 = (n111_tree_20&n110_tree_20)|n109_tree_20;
    assign n110_tree_20 = a_in[10]|b_in[10];

    assign n109_tree_20 = a_in[10]&b_in[10];
    assign n111_tree_20 = (n114_tree_20&n113_tree_20)|n112_tree_20;
    assign n113_tree_20 = a_in[9]|b_in[9];

    assign n112_tree_20 = a_in[9]&b_in[9];
    assign n114_tree_20 = (n117_tree_20&n116_tree_20)|n115_tree_20;
    assign n116_tree_20 = a_in[8]|b_in[8];

    assign n115_tree_20 = a_in[8]&b_in[8];
    assign n117_tree_20 = (n120_tree_20&n119_tree_20)|n118_tree_20;
    assign n119_tree_20 = a_in[7]|b_in[7];

    assign n118_tree_20 = a_in[7]&b_in[7];
    assign n120_tree_20 = (n123_tree_20&n122_tree_20)|n121_tree_20;
    assign n122_tree_20 = a_in[6]|b_in[6];

    assign n121_tree_20 = a_in[6]&b_in[6];
    assign n123_tree_20 = (n126_tree_20&n125_tree_20)|n124_tree_20;
    assign n125_tree_20 = a_in[5]|b_in[5];

    assign n124_tree_20 = a_in[5]&b_in[5];
    assign n126_tree_20 = (n129_tree_20&n128_tree_20)|n127_tree_20;
    assign n128_tree_20 = a_in[4]|b_in[4];

    assign n127_tree_20 = a_in[4]&b_in[4];
    assign n129_tree_20 = (n132_tree_20&n131_tree_20)|n130_tree_20;
    assign n131_tree_20 = a_in[3]|b_in[3];

    assign n130_tree_20 = a_in[3]&b_in[3];
    assign n132_tree_20 = (n135_tree_20&n134_tree_20)|n133_tree_20;
    assign n134_tree_20 = a_in[2]|b_in[2];

    assign n133_tree_20 = a_in[2]&b_in[2];
    assign n135_tree_20 = (n138_tree_20&n137_tree_20)|n136_tree_20;
    assign n137_tree_20 = a_in[1]|b_in[1];

    assign n136_tree_20 = a_in[1]&b_in[1];
    assign n138_tree_20 = a_in[0]&b_in[0];

// adder_forest tree_19
	wire n76_tree_19, n77_tree_19, n78_tree_19, n79_tree_19, n80_tree_19, n81_tree_19, n82_tree_19, n83_tree_19, n84_tree_19, n85_tree_19, n86_tree_19, n87_tree_19, n88_tree_19, n89_tree_19, n90_tree_19, n91_tree_19, n92_tree_19, n93_tree_19, n94_tree_19, n95_tree_19, n96_tree_19, n97_tree_19, n98_tree_19, n99_tree_19, n100_tree_19, n101_tree_19, n102_tree_19, n103_tree_19, n104_tree_19, n105_tree_19, n106_tree_19, n107_tree_19, n108_tree_19, n109_tree_19, n110_tree_19, n111_tree_19, n112_tree_19, n113_tree_19, n114_tree_19, n115_tree_19, n116_tree_19, n117_tree_19, n118_tree_19, n119_tree_19, n120_tree_19, n121_tree_19, n122_tree_19, n123_tree_19, n124_tree_19, n125_tree_19, n126_tree_19, n127_tree_19, n128_tree_19, n129_tree_19, n130_tree_19, n131_tree_19;
    assign sum[19] = n77_tree_19^n76_tree_19;
    assign n76_tree_19 = a_in[19]^b_in[19];
    assign n77_tree_19 = (n80_tree_19&n79_tree_19)|n78_tree_19;
    assign n79_tree_19 = a_in[18]|b_in[18];

    assign n78_tree_19 = a_in[18]&b_in[18];
    assign n80_tree_19 = (n83_tree_19&n82_tree_19)|n81_tree_19;
    assign n82_tree_19 = a_in[17]|b_in[17];

    assign n81_tree_19 = a_in[17]&b_in[17];
    assign n83_tree_19 = (n86_tree_19&n85_tree_19)|n84_tree_19;
    assign n85_tree_19 = a_in[16]|b_in[16];

    assign n84_tree_19 = a_in[16]&b_in[16];
    assign n86_tree_19 = (n89_tree_19&n88_tree_19)|n87_tree_19;
    assign n88_tree_19 = a_in[15]|b_in[15];

    assign n87_tree_19 = a_in[15]&b_in[15];
    assign n89_tree_19 = (n92_tree_19&n91_tree_19)|n90_tree_19;
    assign n91_tree_19 = a_in[14]|b_in[14];

    assign n90_tree_19 = a_in[14]&b_in[14];
    assign n92_tree_19 = (n95_tree_19&n94_tree_19)|n93_tree_19;
    assign n94_tree_19 = a_in[13]|b_in[13];

    assign n93_tree_19 = a_in[13]&b_in[13];
    assign n95_tree_19 = (n98_tree_19&n97_tree_19)|n96_tree_19;
    assign n97_tree_19 = a_in[12]|b_in[12];

    assign n96_tree_19 = a_in[12]&b_in[12];
    assign n98_tree_19 = (n101_tree_19&n100_tree_19)|n99_tree_19;
    assign n100_tree_19 = a_in[11]|b_in[11];

    assign n99_tree_19 = a_in[11]&b_in[11];
    assign n101_tree_19 = (n104_tree_19&n103_tree_19)|n102_tree_19;
    assign n103_tree_19 = a_in[10]|b_in[10];

    assign n102_tree_19 = a_in[10]&b_in[10];
    assign n104_tree_19 = (n107_tree_19&n106_tree_19)|n105_tree_19;
    assign n106_tree_19 = a_in[9]|b_in[9];

    assign n105_tree_19 = a_in[9]&b_in[9];
    assign n107_tree_19 = (n110_tree_19&n109_tree_19)|n108_tree_19;
    assign n109_tree_19 = a_in[8]|b_in[8];

    assign n108_tree_19 = a_in[8]&b_in[8];
    assign n110_tree_19 = (n113_tree_19&n112_tree_19)|n111_tree_19;
    assign n112_tree_19 = a_in[7]|b_in[7];

    assign n111_tree_19 = a_in[7]&b_in[7];
    assign n113_tree_19 = (n116_tree_19&n115_tree_19)|n114_tree_19;
    assign n115_tree_19 = a_in[6]|b_in[6];

    assign n114_tree_19 = a_in[6]&b_in[6];
    assign n116_tree_19 = (n119_tree_19&n118_tree_19)|n117_tree_19;
    assign n118_tree_19 = a_in[5]|b_in[5];

    assign n117_tree_19 = a_in[5]&b_in[5];
    assign n119_tree_19 = (n122_tree_19&n121_tree_19)|n120_tree_19;
    assign n121_tree_19 = a_in[4]|b_in[4];

    assign n120_tree_19 = a_in[4]&b_in[4];
    assign n122_tree_19 = (n125_tree_19&n124_tree_19)|n123_tree_19;
    assign n124_tree_19 = a_in[3]|b_in[3];

    assign n123_tree_19 = a_in[3]&b_in[3];
    assign n125_tree_19 = (n128_tree_19&n127_tree_19)|n126_tree_19;
    assign n127_tree_19 = a_in[2]|b_in[2];

    assign n126_tree_19 = a_in[2]&b_in[2];
    assign n128_tree_19 = (n131_tree_19&n130_tree_19)|n129_tree_19;
    assign n130_tree_19 = a_in[1]|b_in[1];

    assign n129_tree_19 = a_in[1]&b_in[1];
    assign n131_tree_19 = a_in[0]&b_in[0];

// adder_forest tree_18
	wire n72_tree_18, n73_tree_18, n74_tree_18, n75_tree_18, n76_tree_18, n77_tree_18, n78_tree_18, n79_tree_18, n80_tree_18, n81_tree_18, n82_tree_18, n83_tree_18, n84_tree_18, n85_tree_18, n86_tree_18, n87_tree_18, n88_tree_18, n89_tree_18, n90_tree_18, n91_tree_18, n92_tree_18, n93_tree_18, n94_tree_18, n95_tree_18, n96_tree_18, n97_tree_18, n98_tree_18, n99_tree_18, n100_tree_18, n101_tree_18, n102_tree_18, n103_tree_18, n104_tree_18, n105_tree_18, n106_tree_18, n107_tree_18, n108_tree_18, n109_tree_18, n110_tree_18, n111_tree_18, n112_tree_18, n113_tree_18, n114_tree_18, n115_tree_18, n116_tree_18, n117_tree_18, n118_tree_18, n119_tree_18, n120_tree_18, n121_tree_18, n122_tree_18, n123_tree_18, n124_tree_18;
    assign sum[18] = n73_tree_18^n72_tree_18;
    assign n72_tree_18 = a_in[18]^b_in[18];
    assign n73_tree_18 = (n76_tree_18&n75_tree_18)|n74_tree_18;
    assign n75_tree_18 = a_in[17]|b_in[17];

    assign n74_tree_18 = a_in[17]&b_in[17];
    assign n76_tree_18 = (n79_tree_18&n78_tree_18)|n77_tree_18;
    assign n78_tree_18 = a_in[16]|b_in[16];

    assign n77_tree_18 = a_in[16]&b_in[16];
    assign n79_tree_18 = (n82_tree_18&n81_tree_18)|n80_tree_18;
    assign n81_tree_18 = a_in[15]|b_in[15];

    assign n80_tree_18 = a_in[15]&b_in[15];
    assign n82_tree_18 = (n85_tree_18&n84_tree_18)|n83_tree_18;
    assign n84_tree_18 = a_in[14]|b_in[14];

    assign n83_tree_18 = a_in[14]&b_in[14];
    assign n85_tree_18 = (n88_tree_18&n87_tree_18)|n86_tree_18;
    assign n87_tree_18 = a_in[13]|b_in[13];

    assign n86_tree_18 = a_in[13]&b_in[13];
    assign n88_tree_18 = (n91_tree_18&n90_tree_18)|n89_tree_18;
    assign n90_tree_18 = a_in[12]|b_in[12];

    assign n89_tree_18 = a_in[12]&b_in[12];
    assign n91_tree_18 = (n94_tree_18&n93_tree_18)|n92_tree_18;
    assign n93_tree_18 = a_in[11]|b_in[11];

    assign n92_tree_18 = a_in[11]&b_in[11];
    assign n94_tree_18 = (n97_tree_18&n96_tree_18)|n95_tree_18;
    assign n96_tree_18 = a_in[10]|b_in[10];

    assign n95_tree_18 = a_in[10]&b_in[10];
    assign n97_tree_18 = (n100_tree_18&n99_tree_18)|n98_tree_18;
    assign n99_tree_18 = a_in[9]|b_in[9];

    assign n98_tree_18 = a_in[9]&b_in[9];
    assign n100_tree_18 = (n103_tree_18&n102_tree_18)|n101_tree_18;
    assign n102_tree_18 = a_in[8]|b_in[8];

    assign n101_tree_18 = a_in[8]&b_in[8];
    assign n103_tree_18 = (n106_tree_18&n105_tree_18)|n104_tree_18;
    assign n105_tree_18 = a_in[7]|b_in[7];

    assign n104_tree_18 = a_in[7]&b_in[7];
    assign n106_tree_18 = (n109_tree_18&n108_tree_18)|n107_tree_18;
    assign n108_tree_18 = a_in[6]|b_in[6];

    assign n107_tree_18 = a_in[6]&b_in[6];
    assign n109_tree_18 = (n112_tree_18&n111_tree_18)|n110_tree_18;
    assign n111_tree_18 = a_in[5]|b_in[5];

    assign n110_tree_18 = a_in[5]&b_in[5];
    assign n112_tree_18 = (n115_tree_18&n114_tree_18)|n113_tree_18;
    assign n114_tree_18 = a_in[4]|b_in[4];

    assign n113_tree_18 = a_in[4]&b_in[4];
    assign n115_tree_18 = (n118_tree_18&n117_tree_18)|n116_tree_18;
    assign n117_tree_18 = a_in[3]|b_in[3];

    assign n116_tree_18 = a_in[3]&b_in[3];
    assign n118_tree_18 = (n121_tree_18&n120_tree_18)|n119_tree_18;
    assign n120_tree_18 = a_in[2]|b_in[2];

    assign n119_tree_18 = a_in[2]&b_in[2];
    assign n121_tree_18 = (n124_tree_18&n123_tree_18)|n122_tree_18;
    assign n123_tree_18 = a_in[1]|b_in[1];

    assign n122_tree_18 = a_in[1]&b_in[1];
    assign n124_tree_18 = a_in[0]&b_in[0];

// adder_forest tree_17
	wire n68_tree_17, n69_tree_17, n70_tree_17, n71_tree_17, n72_tree_17, n73_tree_17, n74_tree_17, n75_tree_17, n76_tree_17, n77_tree_17, n78_tree_17, n79_tree_17, n80_tree_17, n81_tree_17, n82_tree_17, n83_tree_17, n84_tree_17, n85_tree_17, n86_tree_17, n87_tree_17, n88_tree_17, n89_tree_17, n90_tree_17, n91_tree_17, n92_tree_17, n93_tree_17, n94_tree_17, n95_tree_17, n96_tree_17, n97_tree_17, n98_tree_17, n99_tree_17, n100_tree_17, n101_tree_17, n102_tree_17, n103_tree_17, n104_tree_17, n105_tree_17, n106_tree_17, n107_tree_17, n108_tree_17, n109_tree_17, n110_tree_17, n111_tree_17, n112_tree_17, n113_tree_17, n114_tree_17, n115_tree_17, n116_tree_17, n117_tree_17;
    assign sum[17] = n69_tree_17^n68_tree_17;
    assign n68_tree_17 = a_in[17]^b_in[17];
    assign n69_tree_17 = (n72_tree_17&n71_tree_17)|n70_tree_17;
    assign n71_tree_17 = a_in[16]|b_in[16];

    assign n70_tree_17 = a_in[16]&b_in[16];
    assign n72_tree_17 = (n75_tree_17&n74_tree_17)|n73_tree_17;
    assign n74_tree_17 = a_in[15]|b_in[15];

    assign n73_tree_17 = a_in[15]&b_in[15];
    assign n75_tree_17 = (n78_tree_17&n77_tree_17)|n76_tree_17;
    assign n77_tree_17 = a_in[14]|b_in[14];

    assign n76_tree_17 = a_in[14]&b_in[14];
    assign n78_tree_17 = (n81_tree_17&n80_tree_17)|n79_tree_17;
    assign n80_tree_17 = a_in[13]|b_in[13];

    assign n79_tree_17 = a_in[13]&b_in[13];
    assign n81_tree_17 = (n84_tree_17&n83_tree_17)|n82_tree_17;
    assign n83_tree_17 = a_in[12]|b_in[12];

    assign n82_tree_17 = a_in[12]&b_in[12];
    assign n84_tree_17 = (n87_tree_17&n86_tree_17)|n85_tree_17;
    assign n86_tree_17 = a_in[11]|b_in[11];

    assign n85_tree_17 = a_in[11]&b_in[11];
    assign n87_tree_17 = (n90_tree_17&n89_tree_17)|n88_tree_17;
    assign n89_tree_17 = a_in[10]|b_in[10];

    assign n88_tree_17 = a_in[10]&b_in[10];
    assign n90_tree_17 = (n93_tree_17&n92_tree_17)|n91_tree_17;
    assign n92_tree_17 = a_in[9]|b_in[9];

    assign n91_tree_17 = a_in[9]&b_in[9];
    assign n93_tree_17 = (n96_tree_17&n95_tree_17)|n94_tree_17;
    assign n95_tree_17 = a_in[8]|b_in[8];

    assign n94_tree_17 = a_in[8]&b_in[8];
    assign n96_tree_17 = (n99_tree_17&n98_tree_17)|n97_tree_17;
    assign n98_tree_17 = a_in[7]|b_in[7];

    assign n97_tree_17 = a_in[7]&b_in[7];
    assign n99_tree_17 = (n102_tree_17&n101_tree_17)|n100_tree_17;
    assign n101_tree_17 = a_in[6]|b_in[6];

    assign n100_tree_17 = a_in[6]&b_in[6];
    assign n102_tree_17 = (n105_tree_17&n104_tree_17)|n103_tree_17;
    assign n104_tree_17 = a_in[5]|b_in[5];

    assign n103_tree_17 = a_in[5]&b_in[5];
    assign n105_tree_17 = (n108_tree_17&n107_tree_17)|n106_tree_17;
    assign n107_tree_17 = a_in[4]|b_in[4];

    assign n106_tree_17 = a_in[4]&b_in[4];
    assign n108_tree_17 = (n111_tree_17&n110_tree_17)|n109_tree_17;
    assign n110_tree_17 = a_in[3]|b_in[3];

    assign n109_tree_17 = a_in[3]&b_in[3];
    assign n111_tree_17 = (n114_tree_17&n113_tree_17)|n112_tree_17;
    assign n113_tree_17 = a_in[2]|b_in[2];

    assign n112_tree_17 = a_in[2]&b_in[2];
    assign n114_tree_17 = (n117_tree_17&n116_tree_17)|n115_tree_17;
    assign n116_tree_17 = a_in[1]|b_in[1];

    assign n115_tree_17 = a_in[1]&b_in[1];
    assign n117_tree_17 = a_in[0]&b_in[0];

// adder_forest tree_16
	wire n64_tree_16, n65_tree_16, n66_tree_16, n67_tree_16, n68_tree_16, n69_tree_16, n70_tree_16, n71_tree_16, n72_tree_16, n73_tree_16, n74_tree_16, n75_tree_16, n76_tree_16, n77_tree_16, n78_tree_16, n79_tree_16, n80_tree_16, n81_tree_16, n82_tree_16, n83_tree_16, n84_tree_16, n85_tree_16, n86_tree_16, n87_tree_16, n88_tree_16, n89_tree_16, n90_tree_16, n91_tree_16, n92_tree_16, n93_tree_16, n94_tree_16, n95_tree_16, n96_tree_16, n97_tree_16, n98_tree_16, n99_tree_16, n100_tree_16, n101_tree_16, n102_tree_16, n103_tree_16, n104_tree_16, n105_tree_16, n106_tree_16, n107_tree_16, n108_tree_16, n109_tree_16, n110_tree_16;
    assign sum[16] = n65_tree_16^n64_tree_16;
    assign n64_tree_16 = a_in[16]^b_in[16];
    assign n65_tree_16 = (n68_tree_16&n67_tree_16)|n66_tree_16;
    assign n67_tree_16 = a_in[15]|b_in[15];

    assign n66_tree_16 = a_in[15]&b_in[15];
    assign n68_tree_16 = (n71_tree_16&n70_tree_16)|n69_tree_16;
    assign n70_tree_16 = a_in[14]|b_in[14];

    assign n69_tree_16 = a_in[14]&b_in[14];
    assign n71_tree_16 = (n74_tree_16&n73_tree_16)|n72_tree_16;
    assign n73_tree_16 = a_in[13]|b_in[13];

    assign n72_tree_16 = a_in[13]&b_in[13];
    assign n74_tree_16 = (n77_tree_16&n76_tree_16)|n75_tree_16;
    assign n76_tree_16 = a_in[12]|b_in[12];

    assign n75_tree_16 = a_in[12]&b_in[12];
    assign n77_tree_16 = (n80_tree_16&n79_tree_16)|n78_tree_16;
    assign n79_tree_16 = a_in[11]|b_in[11];

    assign n78_tree_16 = a_in[11]&b_in[11];
    assign n80_tree_16 = (n83_tree_16&n82_tree_16)|n81_tree_16;
    assign n82_tree_16 = a_in[10]|b_in[10];

    assign n81_tree_16 = a_in[10]&b_in[10];
    assign n83_tree_16 = (n86_tree_16&n85_tree_16)|n84_tree_16;
    assign n85_tree_16 = a_in[9]|b_in[9];

    assign n84_tree_16 = a_in[9]&b_in[9];
    assign n86_tree_16 = (n89_tree_16&n88_tree_16)|n87_tree_16;
    assign n88_tree_16 = a_in[8]|b_in[8];

    assign n87_tree_16 = a_in[8]&b_in[8];
    assign n89_tree_16 = (n92_tree_16&n91_tree_16)|n90_tree_16;
    assign n91_tree_16 = a_in[7]|b_in[7];

    assign n90_tree_16 = a_in[7]&b_in[7];
    assign n92_tree_16 = (n95_tree_16&n94_tree_16)|n93_tree_16;
    assign n94_tree_16 = a_in[6]|b_in[6];

    assign n93_tree_16 = a_in[6]&b_in[6];
    assign n95_tree_16 = (n98_tree_16&n97_tree_16)|n96_tree_16;
    assign n97_tree_16 = a_in[5]|b_in[5];

    assign n96_tree_16 = a_in[5]&b_in[5];
    assign n98_tree_16 = (n101_tree_16&n100_tree_16)|n99_tree_16;
    assign n100_tree_16 = a_in[4]|b_in[4];

    assign n99_tree_16 = a_in[4]&b_in[4];
    assign n101_tree_16 = (n104_tree_16&n103_tree_16)|n102_tree_16;
    assign n103_tree_16 = a_in[3]|b_in[3];

    assign n102_tree_16 = a_in[3]&b_in[3];
    assign n104_tree_16 = (n107_tree_16&n106_tree_16)|n105_tree_16;
    assign n106_tree_16 = a_in[2]|b_in[2];

    assign n105_tree_16 = a_in[2]&b_in[2];
    assign n107_tree_16 = (n110_tree_16&n109_tree_16)|n108_tree_16;
    assign n109_tree_16 = a_in[1]|b_in[1];

    assign n108_tree_16 = a_in[1]&b_in[1];
    assign n110_tree_16 = a_in[0]&b_in[0];

// adder_forest tree_15
	wire n60_tree_15, n61_tree_15, n62_tree_15, n63_tree_15, n64_tree_15, n65_tree_15, n66_tree_15, n67_tree_15, n68_tree_15, n69_tree_15, n70_tree_15, n71_tree_15, n72_tree_15, n73_tree_15, n74_tree_15, n75_tree_15, n76_tree_15, n77_tree_15, n78_tree_15, n79_tree_15, n80_tree_15, n81_tree_15, n82_tree_15, n83_tree_15, n84_tree_15, n85_tree_15, n86_tree_15, n87_tree_15, n88_tree_15, n89_tree_15, n90_tree_15, n91_tree_15, n92_tree_15, n93_tree_15, n94_tree_15, n95_tree_15, n96_tree_15, n97_tree_15, n98_tree_15, n99_tree_15, n100_tree_15, n101_tree_15, n102_tree_15, n103_tree_15;
    assign sum[15] = n61_tree_15^n60_tree_15;
    assign n60_tree_15 = a_in[15]^b_in[15];
    assign n61_tree_15 = (n64_tree_15&n63_tree_15)|n62_tree_15;
    assign n63_tree_15 = a_in[14]|b_in[14];

    assign n62_tree_15 = a_in[14]&b_in[14];
    assign n64_tree_15 = (n67_tree_15&n66_tree_15)|n65_tree_15;
    assign n66_tree_15 = a_in[13]|b_in[13];

    assign n65_tree_15 = a_in[13]&b_in[13];
    assign n67_tree_15 = (n70_tree_15&n69_tree_15)|n68_tree_15;
    assign n69_tree_15 = a_in[12]|b_in[12];

    assign n68_tree_15 = a_in[12]&b_in[12];
    assign n70_tree_15 = (n73_tree_15&n72_tree_15)|n71_tree_15;
    assign n72_tree_15 = a_in[11]|b_in[11];

    assign n71_tree_15 = a_in[11]&b_in[11];
    assign n73_tree_15 = (n76_tree_15&n75_tree_15)|n74_tree_15;
    assign n75_tree_15 = a_in[10]|b_in[10];

    assign n74_tree_15 = a_in[10]&b_in[10];
    assign n76_tree_15 = (n79_tree_15&n78_tree_15)|n77_tree_15;
    assign n78_tree_15 = a_in[9]|b_in[9];

    assign n77_tree_15 = a_in[9]&b_in[9];
    assign n79_tree_15 = (n82_tree_15&n81_tree_15)|n80_tree_15;
    assign n81_tree_15 = a_in[8]|b_in[8];

    assign n80_tree_15 = a_in[8]&b_in[8];
    assign n82_tree_15 = (n85_tree_15&n84_tree_15)|n83_tree_15;
    assign n84_tree_15 = a_in[7]|b_in[7];

    assign n83_tree_15 = a_in[7]&b_in[7];
    assign n85_tree_15 = (n88_tree_15&n87_tree_15)|n86_tree_15;
    assign n87_tree_15 = a_in[6]|b_in[6];

    assign n86_tree_15 = a_in[6]&b_in[6];
    assign n88_tree_15 = (n91_tree_15&n90_tree_15)|n89_tree_15;
    assign n90_tree_15 = a_in[5]|b_in[5];

    assign n89_tree_15 = a_in[5]&b_in[5];
    assign n91_tree_15 = (n94_tree_15&n93_tree_15)|n92_tree_15;
    assign n93_tree_15 = a_in[4]|b_in[4];

    assign n92_tree_15 = a_in[4]&b_in[4];
    assign n94_tree_15 = (n97_tree_15&n96_tree_15)|n95_tree_15;
    assign n96_tree_15 = a_in[3]|b_in[3];

    assign n95_tree_15 = a_in[3]&b_in[3];
    assign n97_tree_15 = (n100_tree_15&n99_tree_15)|n98_tree_15;
    assign n99_tree_15 = a_in[2]|b_in[2];

    assign n98_tree_15 = a_in[2]&b_in[2];
    assign n100_tree_15 = (n103_tree_15&n102_tree_15)|n101_tree_15;
    assign n102_tree_15 = a_in[1]|b_in[1];

    assign n101_tree_15 = a_in[1]&b_in[1];
    assign n103_tree_15 = a_in[0]&b_in[0];

// adder_forest tree_14
	wire n56_tree_14, n57_tree_14, n58_tree_14, n59_tree_14, n60_tree_14, n61_tree_14, n62_tree_14, n63_tree_14, n64_tree_14, n65_tree_14, n66_tree_14, n67_tree_14, n68_tree_14, n69_tree_14, n70_tree_14, n71_tree_14, n72_tree_14, n73_tree_14, n74_tree_14, n75_tree_14, n76_tree_14, n77_tree_14, n78_tree_14, n79_tree_14, n80_tree_14, n81_tree_14, n82_tree_14, n83_tree_14, n84_tree_14, n85_tree_14, n86_tree_14, n87_tree_14, n88_tree_14, n89_tree_14, n90_tree_14, n91_tree_14, n92_tree_14, n93_tree_14, n94_tree_14, n95_tree_14, n96_tree_14;
    assign sum[14] = n57_tree_14^n56_tree_14;
    assign n56_tree_14 = a_in[14]^b_in[14];
    assign n57_tree_14 = (n60_tree_14&n59_tree_14)|n58_tree_14;
    assign n59_tree_14 = a_in[13]|b_in[13];

    assign n58_tree_14 = a_in[13]&b_in[13];
    assign n60_tree_14 = (n63_tree_14&n62_tree_14)|n61_tree_14;
    assign n62_tree_14 = a_in[12]|b_in[12];

    assign n61_tree_14 = a_in[12]&b_in[12];
    assign n63_tree_14 = (n66_tree_14&n65_tree_14)|n64_tree_14;
    assign n65_tree_14 = a_in[11]|b_in[11];

    assign n64_tree_14 = a_in[11]&b_in[11];
    assign n66_tree_14 = (n69_tree_14&n68_tree_14)|n67_tree_14;
    assign n68_tree_14 = a_in[10]|b_in[10];

    assign n67_tree_14 = a_in[10]&b_in[10];
    assign n69_tree_14 = (n72_tree_14&n71_tree_14)|n70_tree_14;
    assign n71_tree_14 = a_in[9]|b_in[9];

    assign n70_tree_14 = a_in[9]&b_in[9];
    assign n72_tree_14 = (n75_tree_14&n74_tree_14)|n73_tree_14;
    assign n74_tree_14 = a_in[8]|b_in[8];

    assign n73_tree_14 = a_in[8]&b_in[8];
    assign n75_tree_14 = (n78_tree_14&n77_tree_14)|n76_tree_14;
    assign n77_tree_14 = a_in[7]|b_in[7];

    assign n76_tree_14 = a_in[7]&b_in[7];
    assign n78_tree_14 = (n81_tree_14&n80_tree_14)|n79_tree_14;
    assign n80_tree_14 = a_in[6]|b_in[6];

    assign n79_tree_14 = a_in[6]&b_in[6];
    assign n81_tree_14 = (n84_tree_14&n83_tree_14)|n82_tree_14;
    assign n83_tree_14 = a_in[5]|b_in[5];

    assign n82_tree_14 = a_in[5]&b_in[5];
    assign n84_tree_14 = (n87_tree_14&n86_tree_14)|n85_tree_14;
    assign n86_tree_14 = a_in[4]|b_in[4];

    assign n85_tree_14 = a_in[4]&b_in[4];
    assign n87_tree_14 = (n90_tree_14&n89_tree_14)|n88_tree_14;
    assign n89_tree_14 = a_in[3]|b_in[3];

    assign n88_tree_14 = a_in[3]&b_in[3];
    assign n90_tree_14 = (n93_tree_14&n92_tree_14)|n91_tree_14;
    assign n92_tree_14 = a_in[2]|b_in[2];

    assign n91_tree_14 = a_in[2]&b_in[2];
    assign n93_tree_14 = (n96_tree_14&n95_tree_14)|n94_tree_14;
    assign n95_tree_14 = a_in[1]|b_in[1];

    assign n94_tree_14 = a_in[1]&b_in[1];
    assign n96_tree_14 = a_in[0]&b_in[0];

// adder_forest tree_13
	wire n52_tree_13, n53_tree_13, n54_tree_13, n55_tree_13, n56_tree_13, n57_tree_13, n58_tree_13, n59_tree_13, n60_tree_13, n61_tree_13, n62_tree_13, n63_tree_13, n64_tree_13, n65_tree_13, n66_tree_13, n67_tree_13, n68_tree_13, n69_tree_13, n70_tree_13, n71_tree_13, n72_tree_13, n73_tree_13, n74_tree_13, n75_tree_13, n76_tree_13, n77_tree_13, n78_tree_13, n79_tree_13, n80_tree_13, n81_tree_13, n82_tree_13, n83_tree_13, n84_tree_13, n85_tree_13, n86_tree_13, n87_tree_13, n88_tree_13, n89_tree_13;
    assign sum[13] = n53_tree_13^n52_tree_13;
    assign n52_tree_13 = a_in[13]^b_in[13];
    assign n53_tree_13 = (n56_tree_13&n55_tree_13)|n54_tree_13;
    assign n55_tree_13 = a_in[12]|b_in[12];

    assign n54_tree_13 = a_in[12]&b_in[12];
    assign n56_tree_13 = (n59_tree_13&n58_tree_13)|n57_tree_13;
    assign n58_tree_13 = a_in[11]|b_in[11];

    assign n57_tree_13 = a_in[11]&b_in[11];
    assign n59_tree_13 = (n62_tree_13&n61_tree_13)|n60_tree_13;
    assign n61_tree_13 = a_in[10]|b_in[10];

    assign n60_tree_13 = a_in[10]&b_in[10];
    assign n62_tree_13 = (n65_tree_13&n64_tree_13)|n63_tree_13;
    assign n64_tree_13 = a_in[9]|b_in[9];

    assign n63_tree_13 = a_in[9]&b_in[9];
    assign n65_tree_13 = (n68_tree_13&n67_tree_13)|n66_tree_13;
    assign n67_tree_13 = a_in[8]|b_in[8];

    assign n66_tree_13 = a_in[8]&b_in[8];
    assign n68_tree_13 = (n71_tree_13&n70_tree_13)|n69_tree_13;
    assign n70_tree_13 = a_in[7]|b_in[7];

    assign n69_tree_13 = a_in[7]&b_in[7];
    assign n71_tree_13 = (n74_tree_13&n73_tree_13)|n72_tree_13;
    assign n73_tree_13 = a_in[6]|b_in[6];

    assign n72_tree_13 = a_in[6]&b_in[6];
    assign n74_tree_13 = (n77_tree_13&n76_tree_13)|n75_tree_13;
    assign n76_tree_13 = a_in[5]|b_in[5];

    assign n75_tree_13 = a_in[5]&b_in[5];
    assign n77_tree_13 = (n80_tree_13&n79_tree_13)|n78_tree_13;
    assign n79_tree_13 = a_in[4]|b_in[4];

    assign n78_tree_13 = a_in[4]&b_in[4];
    assign n80_tree_13 = (n83_tree_13&n82_tree_13)|n81_tree_13;
    assign n82_tree_13 = a_in[3]|b_in[3];

    assign n81_tree_13 = a_in[3]&b_in[3];
    assign n83_tree_13 = (n86_tree_13&n85_tree_13)|n84_tree_13;
    assign n85_tree_13 = a_in[2]|b_in[2];

    assign n84_tree_13 = a_in[2]&b_in[2];
    assign n86_tree_13 = (n89_tree_13&n88_tree_13)|n87_tree_13;
    assign n88_tree_13 = a_in[1]|b_in[1];

    assign n87_tree_13 = a_in[1]&b_in[1];
    assign n89_tree_13 = a_in[0]&b_in[0];

// adder_forest tree_12
	wire n48_tree_12, n49_tree_12, n50_tree_12, n51_tree_12, n52_tree_12, n53_tree_12, n54_tree_12, n55_tree_12, n56_tree_12, n57_tree_12, n58_tree_12, n59_tree_12, n60_tree_12, n61_tree_12, n62_tree_12, n63_tree_12, n64_tree_12, n65_tree_12, n66_tree_12, n67_tree_12, n68_tree_12, n69_tree_12, n70_tree_12, n71_tree_12, n72_tree_12, n73_tree_12, n74_tree_12, n75_tree_12, n76_tree_12, n77_tree_12, n78_tree_12, n79_tree_12, n80_tree_12, n81_tree_12, n82_tree_12;
    assign sum[12] = n49_tree_12^n48_tree_12;
    assign n48_tree_12 = a_in[12]^b_in[12];
    assign n49_tree_12 = (n52_tree_12&n51_tree_12)|n50_tree_12;
    assign n51_tree_12 = a_in[11]|b_in[11];

    assign n50_tree_12 = a_in[11]&b_in[11];
    assign n52_tree_12 = (n55_tree_12&n54_tree_12)|n53_tree_12;
    assign n54_tree_12 = a_in[10]|b_in[10];

    assign n53_tree_12 = a_in[10]&b_in[10];
    assign n55_tree_12 = (n58_tree_12&n57_tree_12)|n56_tree_12;
    assign n57_tree_12 = a_in[9]|b_in[9];

    assign n56_tree_12 = a_in[9]&b_in[9];
    assign n58_tree_12 = (n61_tree_12&n60_tree_12)|n59_tree_12;
    assign n60_tree_12 = a_in[8]|b_in[8];

    assign n59_tree_12 = a_in[8]&b_in[8];
    assign n61_tree_12 = (n64_tree_12&n63_tree_12)|n62_tree_12;
    assign n63_tree_12 = a_in[7]|b_in[7];

    assign n62_tree_12 = a_in[7]&b_in[7];
    assign n64_tree_12 = (n67_tree_12&n66_tree_12)|n65_tree_12;
    assign n66_tree_12 = a_in[6]|b_in[6];

    assign n65_tree_12 = a_in[6]&b_in[6];
    assign n67_tree_12 = (n70_tree_12&n69_tree_12)|n68_tree_12;
    assign n69_tree_12 = a_in[5]|b_in[5];

    assign n68_tree_12 = a_in[5]&b_in[5];
    assign n70_tree_12 = (n73_tree_12&n72_tree_12)|n71_tree_12;
    assign n72_tree_12 = a_in[4]|b_in[4];

    assign n71_tree_12 = a_in[4]&b_in[4];
    assign n73_tree_12 = (n76_tree_12&n75_tree_12)|n74_tree_12;
    assign n75_tree_12 = a_in[3]|b_in[3];

    assign n74_tree_12 = a_in[3]&b_in[3];
    assign n76_tree_12 = (n79_tree_12&n78_tree_12)|n77_tree_12;
    assign n78_tree_12 = a_in[2]|b_in[2];

    assign n77_tree_12 = a_in[2]&b_in[2];
    assign n79_tree_12 = (n82_tree_12&n81_tree_12)|n80_tree_12;
    assign n81_tree_12 = a_in[1]|b_in[1];

    assign n80_tree_12 = a_in[1]&b_in[1];
    assign n82_tree_12 = a_in[0]&b_in[0];

// adder_forest tree_11
	wire n44_tree_11, n45_tree_11, n46_tree_11, n47_tree_11, n48_tree_11, n49_tree_11, n50_tree_11, n51_tree_11, n52_tree_11, n53_tree_11, n54_tree_11, n55_tree_11, n56_tree_11, n57_tree_11, n58_tree_11, n59_tree_11, n60_tree_11, n61_tree_11, n62_tree_11, n63_tree_11, n64_tree_11, n65_tree_11, n66_tree_11, n67_tree_11, n68_tree_11, n69_tree_11, n70_tree_11, n71_tree_11, n72_tree_11, n73_tree_11, n74_tree_11, n75_tree_11;
    assign sum[11] = n45_tree_11^n44_tree_11;
    assign n44_tree_11 = a_in[11]^b_in[11];
    assign n45_tree_11 = (n48_tree_11&n47_tree_11)|n46_tree_11;
    assign n47_tree_11 = a_in[10]|b_in[10];

    assign n46_tree_11 = a_in[10]&b_in[10];
    assign n48_tree_11 = (n51_tree_11&n50_tree_11)|n49_tree_11;
    assign n50_tree_11 = a_in[9]|b_in[9];

    assign n49_tree_11 = a_in[9]&b_in[9];
    assign n51_tree_11 = (n54_tree_11&n53_tree_11)|n52_tree_11;
    assign n53_tree_11 = a_in[8]|b_in[8];

    assign n52_tree_11 = a_in[8]&b_in[8];
    assign n54_tree_11 = (n57_tree_11&n56_tree_11)|n55_tree_11;
    assign n56_tree_11 = a_in[7]|b_in[7];

    assign n55_tree_11 = a_in[7]&b_in[7];
    assign n57_tree_11 = (n60_tree_11&n59_tree_11)|n58_tree_11;
    assign n59_tree_11 = a_in[6]|b_in[6];

    assign n58_tree_11 = a_in[6]&b_in[6];
    assign n60_tree_11 = (n63_tree_11&n62_tree_11)|n61_tree_11;
    assign n62_tree_11 = a_in[5]|b_in[5];

    assign n61_tree_11 = a_in[5]&b_in[5];
    assign n63_tree_11 = (n66_tree_11&n65_tree_11)|n64_tree_11;
    assign n65_tree_11 = a_in[4]|b_in[4];

    assign n64_tree_11 = a_in[4]&b_in[4];
    assign n66_tree_11 = (n69_tree_11&n68_tree_11)|n67_tree_11;
    assign n68_tree_11 = a_in[3]|b_in[3];

    assign n67_tree_11 = a_in[3]&b_in[3];
    assign n69_tree_11 = (n72_tree_11&n71_tree_11)|n70_tree_11;
    assign n71_tree_11 = a_in[2]|b_in[2];

    assign n70_tree_11 = a_in[2]&b_in[2];
    assign n72_tree_11 = (n75_tree_11&n74_tree_11)|n73_tree_11;
    assign n74_tree_11 = a_in[1]|b_in[1];

    assign n73_tree_11 = a_in[1]&b_in[1];
    assign n75_tree_11 = a_in[0]&b_in[0];

// adder_forest tree_10
	wire n40_tree_10, n41_tree_10, n42_tree_10, n43_tree_10, n44_tree_10, n45_tree_10, n46_tree_10, n47_tree_10, n48_tree_10, n49_tree_10, n50_tree_10, n51_tree_10, n52_tree_10, n53_tree_10, n54_tree_10, n55_tree_10, n56_tree_10, n57_tree_10, n58_tree_10, n59_tree_10, n60_tree_10, n61_tree_10, n62_tree_10, n63_tree_10, n64_tree_10, n65_tree_10, n66_tree_10, n67_tree_10, n68_tree_10;
    assign sum[10] = n41_tree_10^n40_tree_10;
    assign n40_tree_10 = a_in[10]^b_in[10];
    assign n41_tree_10 = (n44_tree_10&n43_tree_10)|n42_tree_10;
    assign n43_tree_10 = a_in[9]|b_in[9];

    assign n42_tree_10 = a_in[9]&b_in[9];
    assign n44_tree_10 = (n47_tree_10&n46_tree_10)|n45_tree_10;
    assign n46_tree_10 = a_in[8]|b_in[8];

    assign n45_tree_10 = a_in[8]&b_in[8];
    assign n47_tree_10 = (n50_tree_10&n49_tree_10)|n48_tree_10;
    assign n49_tree_10 = a_in[7]|b_in[7];

    assign n48_tree_10 = a_in[7]&b_in[7];
    assign n50_tree_10 = (n53_tree_10&n52_tree_10)|n51_tree_10;
    assign n52_tree_10 = a_in[6]|b_in[6];

    assign n51_tree_10 = a_in[6]&b_in[6];
    assign n53_tree_10 = (n56_tree_10&n55_tree_10)|n54_tree_10;
    assign n55_tree_10 = a_in[5]|b_in[5];

    assign n54_tree_10 = a_in[5]&b_in[5];
    assign n56_tree_10 = (n59_tree_10&n58_tree_10)|n57_tree_10;
    assign n58_tree_10 = a_in[4]|b_in[4];

    assign n57_tree_10 = a_in[4]&b_in[4];
    assign n59_tree_10 = (n62_tree_10&n61_tree_10)|n60_tree_10;
    assign n61_tree_10 = a_in[3]|b_in[3];

    assign n60_tree_10 = a_in[3]&b_in[3];
    assign n62_tree_10 = (n65_tree_10&n64_tree_10)|n63_tree_10;
    assign n64_tree_10 = a_in[2]|b_in[2];

    assign n63_tree_10 = a_in[2]&b_in[2];
    assign n65_tree_10 = (n68_tree_10&n67_tree_10)|n66_tree_10;
    assign n67_tree_10 = a_in[1]|b_in[1];

    assign n66_tree_10 = a_in[1]&b_in[1];
    assign n68_tree_10 = a_in[0]&b_in[0];

// adder_forest tree_9
	wire n36_tree_9, n37_tree_9, n38_tree_9, n39_tree_9, n40_tree_9, n41_tree_9, n42_tree_9, n43_tree_9, n44_tree_9, n45_tree_9, n46_tree_9, n47_tree_9, n48_tree_9, n49_tree_9, n50_tree_9, n51_tree_9, n52_tree_9, n53_tree_9, n54_tree_9, n55_tree_9, n56_tree_9, n57_tree_9, n58_tree_9, n59_tree_9, n60_tree_9, n61_tree_9;
    assign sum[9] = n37_tree_9^n36_tree_9;
    assign n36_tree_9 = a_in[9]^b_in[9];
    assign n37_tree_9 = (n40_tree_9&n39_tree_9)|n38_tree_9;
    assign n39_tree_9 = a_in[8]|b_in[8];

    assign n38_tree_9 = a_in[8]&b_in[8];
    assign n40_tree_9 = (n43_tree_9&n42_tree_9)|n41_tree_9;
    assign n42_tree_9 = a_in[7]|b_in[7];

    assign n41_tree_9 = a_in[7]&b_in[7];
    assign n43_tree_9 = (n46_tree_9&n45_tree_9)|n44_tree_9;
    assign n45_tree_9 = a_in[6]|b_in[6];

    assign n44_tree_9 = a_in[6]&b_in[6];
    assign n46_tree_9 = (n49_tree_9&n48_tree_9)|n47_tree_9;
    assign n48_tree_9 = a_in[5]|b_in[5];

    assign n47_tree_9 = a_in[5]&b_in[5];
    assign n49_tree_9 = (n52_tree_9&n51_tree_9)|n50_tree_9;
    assign n51_tree_9 = a_in[4]|b_in[4];

    assign n50_tree_9 = a_in[4]&b_in[4];
    assign n52_tree_9 = (n55_tree_9&n54_tree_9)|n53_tree_9;
    assign n54_tree_9 = a_in[3]|b_in[3];

    assign n53_tree_9 = a_in[3]&b_in[3];
    assign n55_tree_9 = (n58_tree_9&n57_tree_9)|n56_tree_9;
    assign n57_tree_9 = a_in[2]|b_in[2];

    assign n56_tree_9 = a_in[2]&b_in[2];
    assign n58_tree_9 = (n61_tree_9&n60_tree_9)|n59_tree_9;
    assign n60_tree_9 = a_in[1]|b_in[1];

    assign n59_tree_9 = a_in[1]&b_in[1];
    assign n61_tree_9 = a_in[0]&b_in[0];

// adder_forest tree_8
	wire n32_tree_8, n33_tree_8, n34_tree_8, n35_tree_8, n36_tree_8, n37_tree_8, n38_tree_8, n39_tree_8, n40_tree_8, n41_tree_8, n42_tree_8, n43_tree_8, n44_tree_8, n45_tree_8, n46_tree_8, n47_tree_8, n48_tree_8, n49_tree_8, n50_tree_8, n51_tree_8, n52_tree_8, n53_tree_8, n54_tree_8;
    assign sum[8] = n33_tree_8^n32_tree_8;
    assign n32_tree_8 = a_in[8]^b_in[8];
    assign n33_tree_8 = (n36_tree_8&n35_tree_8)|n34_tree_8;
    assign n35_tree_8 = a_in[7]|b_in[7];

    assign n34_tree_8 = a_in[7]&b_in[7];
    assign n36_tree_8 = (n39_tree_8&n38_tree_8)|n37_tree_8;
    assign n38_tree_8 = a_in[6]|b_in[6];

    assign n37_tree_8 = a_in[6]&b_in[6];
    assign n39_tree_8 = (n42_tree_8&n41_tree_8)|n40_tree_8;
    assign n41_tree_8 = a_in[5]|b_in[5];

    assign n40_tree_8 = a_in[5]&b_in[5];
    assign n42_tree_8 = (n45_tree_8&n44_tree_8)|n43_tree_8;
    assign n44_tree_8 = a_in[4]|b_in[4];

    assign n43_tree_8 = a_in[4]&b_in[4];
    assign n45_tree_8 = (n48_tree_8&n47_tree_8)|n46_tree_8;
    assign n47_tree_8 = a_in[3]|b_in[3];

    assign n46_tree_8 = a_in[3]&b_in[3];
    assign n48_tree_8 = (n51_tree_8&n50_tree_8)|n49_tree_8;
    assign n50_tree_8 = a_in[2]|b_in[2];

    assign n49_tree_8 = a_in[2]&b_in[2];
    assign n51_tree_8 = (n54_tree_8&n53_tree_8)|n52_tree_8;
    assign n53_tree_8 = a_in[1]|b_in[1];

    assign n52_tree_8 = a_in[1]&b_in[1];
    assign n54_tree_8 = a_in[0]&b_in[0];

// adder_forest tree_7
	wire n28_tree_7, n29_tree_7, n30_tree_7, n31_tree_7, n32_tree_7, n33_tree_7, n34_tree_7, n35_tree_7, n36_tree_7, n37_tree_7, n38_tree_7, n39_tree_7, n40_tree_7, n41_tree_7, n42_tree_7, n43_tree_7, n44_tree_7, n45_tree_7, n46_tree_7, n47_tree_7;
    assign sum[7] = n29_tree_7^n28_tree_7;
    assign n28_tree_7 = a_in[7]^b_in[7];
    assign n29_tree_7 = (n32_tree_7&n31_tree_7)|n30_tree_7;
    assign n31_tree_7 = a_in[6]|b_in[6];

    assign n30_tree_7 = a_in[6]&b_in[6];
    assign n32_tree_7 = (n35_tree_7&n34_tree_7)|n33_tree_7;
    assign n34_tree_7 = a_in[5]|b_in[5];

    assign n33_tree_7 = a_in[5]&b_in[5];
    assign n35_tree_7 = (n38_tree_7&n37_tree_7)|n36_tree_7;
    assign n37_tree_7 = a_in[4]|b_in[4];

    assign n36_tree_7 = a_in[4]&b_in[4];
    assign n38_tree_7 = (n41_tree_7&n40_tree_7)|n39_tree_7;
    assign n40_tree_7 = a_in[3]|b_in[3];

    assign n39_tree_7 = a_in[3]&b_in[3];
    assign n41_tree_7 = (n44_tree_7&n43_tree_7)|n42_tree_7;
    assign n43_tree_7 = a_in[2]|b_in[2];

    assign n42_tree_7 = a_in[2]&b_in[2];
    assign n44_tree_7 = (n47_tree_7&n46_tree_7)|n45_tree_7;
    assign n46_tree_7 = a_in[1]|b_in[1];

    assign n45_tree_7 = a_in[1]&b_in[1];
    assign n47_tree_7 = a_in[0]&b_in[0];

// adder_forest tree_6
	wire n24_tree_6, n25_tree_6, n26_tree_6, n27_tree_6, n28_tree_6, n29_tree_6, n30_tree_6, n31_tree_6, n32_tree_6, n33_tree_6, n34_tree_6, n35_tree_6, n36_tree_6, n37_tree_6, n38_tree_6, n39_tree_6, n40_tree_6;
    assign sum[6] = n25_tree_6^n24_tree_6;
    assign n24_tree_6 = a_in[6]^b_in[6];
    assign n25_tree_6 = (n28_tree_6&n27_tree_6)|n26_tree_6;
    assign n27_tree_6 = a_in[5]|b_in[5];

    assign n26_tree_6 = a_in[5]&b_in[5];
    assign n28_tree_6 = (n31_tree_6&n30_tree_6)|n29_tree_6;
    assign n30_tree_6 = a_in[4]|b_in[4];

    assign n29_tree_6 = a_in[4]&b_in[4];
    assign n31_tree_6 = (n34_tree_6&n33_tree_6)|n32_tree_6;
    assign n33_tree_6 = a_in[3]|b_in[3];

    assign n32_tree_6 = a_in[3]&b_in[3];
    assign n34_tree_6 = (n37_tree_6&n36_tree_6)|n35_tree_6;
    assign n36_tree_6 = a_in[2]|b_in[2];

    assign n35_tree_6 = a_in[2]&b_in[2];
    assign n37_tree_6 = (n40_tree_6&n39_tree_6)|n38_tree_6;
    assign n39_tree_6 = a_in[1]|b_in[1];

    assign n38_tree_6 = a_in[1]&b_in[1];
    assign n40_tree_6 = a_in[0]&b_in[0];

// adder_forest tree_5
	wire n20_tree_5, n21_tree_5, n22_tree_5, n23_tree_5, n24_tree_5, n25_tree_5, n26_tree_5, n27_tree_5, n28_tree_5, n29_tree_5, n30_tree_5, n31_tree_5, n32_tree_5, n33_tree_5;
    assign sum[5] = n21_tree_5^n20_tree_5;
    assign n20_tree_5 = a_in[5]^b_in[5];
    assign n21_tree_5 = (n24_tree_5&n23_tree_5)|n22_tree_5;
    assign n23_tree_5 = a_in[4]|b_in[4];

    assign n22_tree_5 = a_in[4]&b_in[4];
    assign n24_tree_5 = (n27_tree_5&n26_tree_5)|n25_tree_5;
    assign n26_tree_5 = a_in[3]|b_in[3];

    assign n25_tree_5 = a_in[3]&b_in[3];
    assign n27_tree_5 = (n30_tree_5&n29_tree_5)|n28_tree_5;
    assign n29_tree_5 = a_in[2]|b_in[2];

    assign n28_tree_5 = a_in[2]&b_in[2];
    assign n30_tree_5 = (n33_tree_5&n32_tree_5)|n31_tree_5;
    assign n32_tree_5 = a_in[1]|b_in[1];

    assign n31_tree_5 = a_in[1]&b_in[1];
    assign n33_tree_5 = a_in[0]&b_in[0];

// adder_forest tree_4
	wire n16_tree_4, n17_tree_4, n18_tree_4, n19_tree_4, n20_tree_4, n21_tree_4, n22_tree_4, n23_tree_4, n24_tree_4, n25_tree_4, n26_tree_4;
    assign sum[4] = n17_tree_4^n16_tree_4;
    assign n16_tree_4 = a_in[4]^b_in[4];
    assign n17_tree_4 = (n20_tree_4&n19_tree_4)|n18_tree_4;
    assign n19_tree_4 = a_in[3]|b_in[3];

    assign n18_tree_4 = a_in[3]&b_in[3];
    assign n20_tree_4 = (n23_tree_4&n22_tree_4)|n21_tree_4;
    assign n22_tree_4 = a_in[2]|b_in[2];

    assign n21_tree_4 = a_in[2]&b_in[2];
    assign n23_tree_4 = (n26_tree_4&n25_tree_4)|n24_tree_4;
    assign n25_tree_4 = a_in[1]|b_in[1];

    assign n24_tree_4 = a_in[1]&b_in[1];
    assign n26_tree_4 = a_in[0]&b_in[0];

// adder_forest tree_3
	wire n12_tree_3, n13_tree_3, n14_tree_3, n15_tree_3, n16_tree_3, n17_tree_3, n18_tree_3, n19_tree_3;
    assign sum[3] = n13_tree_3^n12_tree_3;
    assign n12_tree_3 = a_in[3]^b_in[3];
    assign n13_tree_3 = (n16_tree_3&n15_tree_3)|n14_tree_3;
    assign n15_tree_3 = a_in[2]|b_in[2];

    assign n14_tree_3 = a_in[2]&b_in[2];
    assign n16_tree_3 = (n19_tree_3&n18_tree_3)|n17_tree_3;
    assign n18_tree_3 = a_in[1]|b_in[1];

    assign n17_tree_3 = a_in[1]&b_in[1];
    assign n19_tree_3 = a_in[0]&b_in[0];

// adder_forest tree_2
	wire n8_tree_2, n9_tree_2, n10_tree_2, n11_tree_2, n12_tree_2;
    assign sum[2] = n9_tree_2^n8_tree_2;
    assign n8_tree_2 = a_in[2]^b_in[2];
    assign n9_tree_2 = (n12_tree_2&n11_tree_2)|n10_tree_2;
    assign n11_tree_2 = a_in[1]|b_in[1];

    assign n10_tree_2 = a_in[1]&b_in[1];
    assign n12_tree_2 = a_in[0]&b_in[0];

// adder_forest tree_1
	wire n4_tree_1, n5_tree_1;
    assign sum[1] = n5_tree_1^n4_tree_1;
    assign n4_tree_1 = a_in[1]^b_in[1];
    assign n5_tree_1 = a_in[0]&b_in[0];

// adder_forest tree_0
	wire n3_tree_0;
	assign sum[0] = n3_tree_0;
    assign n3_tree_0 = a_in[0]^b_in[0];

endmodule // ripple_carry
