magic
tech sky130A
magscale 1 2
timestamp 1652882935
<< obsli1 >>
rect 1104 2159 8832 7633
<< obsm1 >>
rect 14 2128 8832 7664
<< metal2 >>
rect 1278 9200 1390 10000
rect 7074 9200 7186 10000
rect -10 0 102 800
rect 5142 0 5254 800
<< obsm2 >>
rect 20 9144 1222 9200
rect 1446 9144 7018 9200
rect 7242 9144 8078 9200
rect 20 856 8078 9144
rect 158 711 5086 856
rect 5310 711 8078 856
<< metal3 >>
rect 9200 6748 10000 6988
rect 0 5388 800 5628
rect 9200 628 10000 868
<< obsm3 >>
rect 800 7068 9200 7649
rect 800 6668 9120 7068
rect 800 5708 9200 6668
rect 880 5308 9200 5708
rect 800 948 9200 5308
rect 800 715 9120 948
<< metal4 >>
rect 2242 2128 2562 7664
rect 3542 2128 3862 7664
rect 4840 2128 5160 7664
rect 6139 2128 6459 7664
rect 7437 2128 7757 7664
<< obsm4 >>
rect 3942 2128 4760 7664
rect 5240 2128 6059 7664
<< labels >>
rlabel metal3 s 9200 6748 10000 6988 6 chain
port 1 nsew signal output
rlabel metal2 s 5142 0 5254 800 6 clk
port 2 nsew signal input
rlabel metal3 s 0 5388 800 5628 6 outputs[0]
port 3 nsew signal output
rlabel metal2 s -10 0 102 800 6 outputs[1]
port 4 nsew signal output
rlabel metal2 s 1278 9200 1390 10000 6 outputs[2]
port 5 nsew signal output
rlabel metal2 s 7074 9200 7186 10000 6 outputs[3]
port 6 nsew signal output
rlabel metal3 s 9200 628 10000 868 6 reset
port 7 nsew signal input
rlabel metal4 s 2242 2128 2562 7664 6 vccd1
port 8 nsew power input
rlabel metal4 s 4840 2128 5160 7664 6 vccd1
port 8 nsew power input
rlabel metal4 s 7437 2128 7757 7664 6 vccd1
port 8 nsew power input
rlabel metal4 s 3542 2128 3862 7664 6 vssd1
port 9 nsew ground input
rlabel metal4 s 6139 2128 6459 7664 6 vssd1
port 9 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 10000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 205242
string GDS_FILE /openlane/designs/wrapped_instrumented_adder/runs/RUN_2022.05.18_14.08.09/results/finishing/instrumented_adder.magic.gds
string GDS_START 114290
<< end >>

